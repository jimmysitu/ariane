/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 3561;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd0080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h08090000_38000000,
        64'hda0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'hffffb2c6_ffffb962,
        64'hffffb962_ffffb2c6,
        64'hffffb962_ffffb74c,
        64'hffffb962_ffffb962,
        64'hffffb886_ffffb2c6,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb2c6,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb2c6_ffffb688,
        64'hffffb2c6_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb2c6_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb962,
        64'hffffb962_ffffb936,
        64'hffffb2b0_ffffb2c8,
        64'hffffb2c8_ffffb2c8,
        64'hffffb2c8_ffffb2c8,
        64'hffffb280_ffffb2c8,
        64'hffffb2c8_ffffb2c8,
        64'hffffb2c8_ffffb2c8,
        64'hffffb2c8_ffffb2c8,
        64'hffffb200_ffffb2c8,
        64'hffffb298_ffffb2c8,
        64'hffffb240_ffffb04c,
        64'hffffb0e2_ffffb0e2,
        64'hffffb06a_ffffb0e2,
        64'hffffb088_ffffb0e2,
        64'hffffb0e2_ffffb0e2,
        64'hffffb0e2_ffffb0e2,
        64'hffffb0e2_ffffb0e2,
        64'hffffb0c4_ffffb0e2,
        64'hffffb0e2_ffffb0a6,
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_0000000a,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00586c6c_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000000_00007525,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000000_00007525,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_58323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h000a5838_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h000a5838_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_000a586c,
        64'h6c363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h00000000_0a756c6c,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h00000000_0a756c6c,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_0a583830,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_0a583830,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_0a583830,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_0a583830,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h000a586c_6c363130,
        64'h25202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h000a5832_3025202c,
        64'h58323025_202c5832,
        64'h3025202c_58323025,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h00000000_0a642520,
        64'h3a737574_61747320,
        64'h2c64656c_69616620,
        64'h64616552_20304453,
        64'h00000000_0a216465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a6425,
        64'h203a7375_74617473,
        64'h202c6465_6c696166,
        64'h206e6f69_74617a69,
        64'h6c616974_696e6920,
        64'h64726163_20304453,
        64'h0000000a_6425203a,
        64'h73757461_7473202c,
        64'h64656c69_6166206c,
        64'h61697469_6e692067,
        64'h69666e6f_63204453,
        64'h00000000_0000000a,
        64'h2164656c_69616620,
        64'h6769666e_6f632070,
        64'h756b6f6f_6c204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000a2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_262394cf,
        64'hc0ef4505_a031fef4,
        64'h26234785_e7892781,
        64'h0807f793_278187aa,
        64'ha31fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'h0001a011_f6e7fee3,
        64'h02700793_0ff7f713,
        64'hfe944783_fef404a3,
        64'h2785fe94_4783cf99,
        64'h27810407_f7932781,
        64'h87aaa6bf_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h3783a0ad_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'ha61fd0ef_fd843503,
        64'h50078593_67854601,
        64'h4685a829_fef42623,
        64'h87aaa7bf_d0effd84,
        64'h35033007_85936785,
        64'h46014685_00f71f63,
        64'h4785873e_0347c783,
        64'hfd843783_a8adfe04,
        64'h04a3a08f_c0ef4505,
        64'hb13fe0ef_853e03e0,
        64'h0593863a_fe645703,
        64'h43dcfd84_3783fef4,
        64'h13230407_e793fe64,
        64'h5783fef4_132387aa,
        64'hb01fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'h86e79523_47411ffe,
        64'hb797b55f_e0ef853e,
        64'h4591863a_fea45703,
        64'h43dcfd84_3783fef4,
        64'h15238ff9_17fd6785,
        64'hfea45703_fef41523,
        64'h0017979b_fea45783,
        64'haa354785_8ae7a123,
        64'h47051ffe_b79787af,
        64'hc0ef8225_05130000,
        64'h151781a5_85930000,
        64'h159748e0_0613a025,
        64'h02f71c63_478d873e,
        64'h0377c783_fd843783,
        64'hfef41523_04000793,
        64'h8c07ae23_1ffeb797,
        64'ha2514785_8ee7a523,
        64'h47051ffe_b7978c2f,
        64'hc0ef86a5_05130000,
        64'h15178625_85930000,
        64'h159748d0_0613a025,
        64'h04f71763_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_9207a023,
        64'h1ffeb797_c385fd84,
        64'h3783fca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'hb8ffe0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_c4ffe0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe842783,
        64'ha83dfef4_26234785,
        64'hc73fe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe84,
        64'h2703fef4_242387aa,
        64'hc61fe0ef_853e0300,
        64'h059343dc_fd843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aac57f,
        64'hd0effd84_35036000,
        64'h0593863e_4681fd44,
        64'h2783fcf4_2a2387ae,
        64'hfca43c23_1800f022,
        64'hf4067179_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aac55f,
        64'he0ef853e_93811782,
        64'h278127c1_43dcfc84,
        64'h3783d15f_e0ef853e,
        64'h03000593_460943dc,
        64'hfc843783_dfc52781,
        64'h8b89fdc4_2783a83d,
        64'hfef42623_4785d39f,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfc843783_c3852781,
        64'h8ff967a1_fdc42703,
        64'hfcf42e23_87aad27f,
        64'he0ef853e_03000593,
        64'h43dcfc84_3783a8bd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_d1dfd0ef,
        64'hfc843503_80078593,
        64'h6785863e_4685fe44,
        64'h2783aae7_9e234745,
        64'h1ffeb797_f56fe0ef,
        64'hfc843503_85befc04,
        64'h36032781_fe245783,
        64'hdbbfe0ef_853e4591,
        64'h863afe04_570343dc,
        64'hfc843783_fef41023,
        64'h8ff917fd_6785fe04,
        64'h5703fef4_10232000,
        64'h0793fef4_11234785,
        64'hfce7dee3_1ff00793,
        64'h0007871b_fe842783,
        64'hfef42423_2785fe84,
        64'h27830007_802397ba,
        64'hfc043703_fe842783,
        64'ha2154785_b2e7a923,
        64'h47051ffe_b797b0af,
        64'hc0efab25_05130000,
        64'h1517aaa5_85930000,
        64'h159735d0_0613a081,
        64'hfe042423_b407ac23,
        64'h1ffeb797_aaa14785,
        64'hb6e7a323_47051ffe,
        64'hb797b3ef_c0efae65,
        64'h05130000_1517ade5,
        64'h85930000_159735c0,
        64'h0613a025_02f71d63,
        64'h11178793_111117b7,
        64'h873e53dc_fc843783,
        64'hb807ae23_1ffeb797,
        64'hc385fc84_3783fe04,
        64'h2223fcb4_3023fca4,
        64'h34230080_f822fc06,
        64'h71398082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_a019fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aae63f_d0effd84,
        64'h3503a007_859367ad,
        64'h46014681_a03dfef4,
        64'h26234785_a82d4785,
        64'hc0e7a323_47051ffe,
        64'hb797bdef_c0efb865,
        64'h05130000_1517b7e5,
        64'h85930000_159732d0,
        64'h0613a025_cb8d2781,
        64'hfec42783_fef42623,
        64'h87aaeb3f_d0effd84,
        64'h35037007_8593678d,
        64'h863e4681_4bbcfd84,
        64'h3783c407_a7231ffe,
        64'hb797a841_4785c4e7,
        64'hae234705_1ffeb797,
        64'hc34fc0ef_bdc50513,
        64'h00001517_bd458593,
        64'h00001597_32c00613,
        64'ha02504f7_1e631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783c807,
        64'ha9231ffe_b797c385,
        64'hfd843783_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efe84_2783fe04,
        64'h2423fa5f_e0ef853a,
        64'h02c00593_863e93c1,
        64'h17c20047_e793fe44,
        64'h578343d8_fd843783,
        64'hfef41223_87aaf8ff,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783d3e5,
        64'h27818b89_2781fe64,
        64'h5783fef4_132387aa,
        64'hfb1fe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'ha821fef4_132387aa,
        64'hfc9fe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'h812ff0ef_853e02c0,
        64'h0593863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12230017_e79393c1,
        64'h17c28fd9_fe445783,
        64'hfec45703_fef41623,
        64'hf007f793_fec45783,
        64'hfef41623_0087979b,
        64'hfec45783_fef41223,
        64'h0ff7f793_fe445783,
        64'hfef41223_87aa82ef,
        64'hf0ef853e_02c00593,
        64'h43dcfd84_3783a0a5,
        64'h87aff0ef_853e02c0,
        64'h0593863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12230017_e79393c1,
        64'h17c28fd9_fe445783,
        64'h93410307_97138fd9,
        64'hfe245783_fec45703,
        64'hfef41623_f007f793,
        64'hfec45783_fef41623,
        64'h0087979b_fec45783,
        64'hfef41123_0c07f793,
        64'hfe245783_fef41123,
        64'h0067979b_fe245783,
        64'hfef41123_0087d79b,
        64'hfec45783_fef41223,
        64'h03f7f793_fe445783,
        64'hfef41223_87aa8c6f,
        64'hf0ef853e_02c00593,
        64'h43dcfd84_378308f7,
        64'h1e634789_873e0367,
        64'hc783fd84_3783a249,
        64'hfef42423_478500e7,
        64'hf6631000_07930007,
        64'h871bfee4_5783fae7,
        64'hfee31000_07930007,
        64'h871bfee4_5783fef4,
        64'h17230017_979bfee4,
        64'h5783a839_fef41623,
        64'h0017d79b_fee45783,
        64'h00e7e963_2781fd44,
        64'h27830007_871b02f7,
        64'h57bb2781_fee45783,
        64'h4798fd84_3783a82d,
        64'hfef41723_4785a2ed,
        64'hfef42423_478506e7,
        64'hfa637fe0_07930007,
        64'h871bfee4_5783fae7,
        64'hffe37fe0_07930007,
        64'h871bfee4_5783fef4,
        64'h17232785_fee45783,
        64'ha831fef4_16230017,
        64'hd79bfee4_578300e7,
        64'he9632781_fd442783,
        64'h0007871b_02f757bb,
        64'h2781fee4_57834798,
        64'hfd843783_a825fef4,
        64'h17234785_ac914785,
        64'hf0e7a723_47051ffe,
        64'hb797ee6f_c0efe8e5,
        64'h05130000_1517e865,
        64'h85930000_15972b80,
        64'h0613a025_08f71963,
        64'h4789873e_0367c783,
        64'hfd843783_a26ff0ef,
        64'h853e02c0_0593863a,
        64'hfe445703_43dcfd84,
        64'h3783fef4_12239be9,
        64'hfe445783_fef41223,
        64'h87aaa12f_f0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783f607_ab231ffe,
        64'hb797a4e9_4785f8e7,
        64'ha2234705_1ffeb797,
        64'hf5cfc0ef_f0450513,
        64'h00001517_efc58593,
        64'h00001597_2b700613,
        64'ha02506f7_1e631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783fa07,
        64'had231ffe_b797c385,
        64'hfd843783_fe041623,
        64'hfcf42a23_87aefca4,
        64'h3c231800_f022f406,
        64'h71798082_61657406,
        64'h70a6853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_a32ff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_f9843783,
        64'hb72ff0ef_853e0280,
        64'h0593863a_0ff77713,
        64'hfe442703_43dcf984,
        64'h3783fef4_22230047,
        64'he793fe44_2783fef4,
        64'h222387aa_b64ff0ef,
        64'h853e0280_059343dc,
        64'hf9843783_a2bfc0ef,
        64'h3e800513_a09dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa7300_00eff984,
        64'h350302f7_1163479d,
        64'h873e57fc_f9843783,
        64'ha849fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa0b80,
        64'h00eff984_350385be,
        64'h5f9cf984_3783b88f,
        64'hf0ef853e_03000593,
        64'h460943dc_f9843783,
        64'hdfc52781_8b89fe44,
        64'h2783a8d1_fef42623,
        64'h4785bacf_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_f9843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aab9af_f0ef853e,
        64'h03000593_43dcf984,
        64'h3783aa11_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hb90fe0ef_f9843503,
        64'h60000593_863e4681,
        64'hfe842783_df985007,
        64'h071b0319_7737f984,
        64'h3783fef4_24231007,
        64'h879b03b9_07b7a831,
        64'hdf985007_071b0319,
        64'h7737f984_3783fef4,
        64'h24231007_879b03b9,
        64'h07b702f7_10634791,
        64'h873e57fc_f9843783,
        64'ha099df98_2007071b,
        64'h0bebc737_f9843783,
        64'hfef42423_2007879b,
        64'h03b907b7_02f71063,
        64'h479d873e_57fcf984,
        64'h3783a275_fef42623,
        64'h47851407_89632781,
        64'hfec42783_fef42623,
        64'h87aa1d40_00eff984,
        64'h35035007_85930319,
        64'h77b7df98_5007071b,
        64'h03197737_f9843783,
        64'hcb2ff0ef_853e0300,
        64'h05934609_43dcf984,
        64'h3783dfc5_27818b89,
        64'hfe442783_aafdfef4,
        64'h26234785_cd6ff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8f984,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_cc4ff0ef,
        64'h853e0300_059343dc,
        64'hf9843783_ac3dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aacbaf_e0eff984,
        64'h35036000_0593863e,
        64'h4681fe84_2783fef4,
        64'h24231007_879b03b9,
        64'h07b70cf7_16634789,
        64'h873e0347_c783f984,
        64'h3783a451_fef42623,
        64'h47852207_85632781,
        64'hfec42783_fef42623,
        64'h87aa2ac0_00eff984,
        64'h350385be_5f9cf984,
        64'h3783df98_0807071b,
        64'h02faf737_f9843783,
        64'hd8aff0ef_853e0300,
        64'h05934609_43dcf984,
        64'h3783dfc5_27818b89,
        64'hfe442783_acd9fef4,
        64'h26234785_daeff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8f984,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_d9cff0ef,
        64'h853e0300_059343dc,
        64'hf9843783_ae19fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aad92f_e0eff984,
        64'h35036000_0593863e,
        64'h4685fe84_2783fef4,
        64'h242337c5_810007b7,
        64'h32e79d23_47451ffe,
        64'hb797fd5f_e0eff984,
        64'h350385be_863afa04,
        64'h07132781_fe245783,
        64'he3aff0ef_853e4591,
        64'h863afe04_570343dc,
        64'hf9843783_fef41023,
        64'h8ff917fd_6785fe04,
        64'h5703fef4_10230400,
        64'h0793fef4_11234785,
        64'hae794785_38e7a523,
        64'h47051ffe_b797b63f,
        64'hc0ef30a5_05130000,
        64'h15173025_85930000,
        64'h15971f40_0613a025,
        64'h14f71163_4785873e,
        64'h0347c783_f9843783,
        64'h3a07ae23_1ffeb797,
        64'haef94785_3ce7a523,
        64'h47051ffe_b797ba3f,
        64'hc0ef34a5_05130000,
        64'h15173425_85930000,
        64'h15971f30_0613a025,
        64'h04f71363_11178793,
        64'h111117b7_873e53dc,
        64'hf9843783_4007a023,
        64'h1ffeb797_c385f984,
        64'h3783fc04_3c23fc04,
        64'h3823fc04_3423fc04,
        64'h3023fa04_3c23fa04,
        64'h3823fa04_3423fa04,
        64'h3023f8a4_3c231880,
        64'hf0a2f486_71598082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'he8eff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfc843783_f4eff0ef,
        64'h853e0300_05934609,
        64'h43dcfc84_3783dfc5,
        64'h27818b89_fdc42783,
        64'ha83dfef4_26234785,
        64'hf72ff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fc84_3783c385,
        64'h27818ff9_67a1fdc4,
        64'h2703fcf4_2e2387aa,
        64'hf60ff0ef_853e0300,
        64'h059343dc_fc843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaf56f,
        64'he0effc84_35036000,
        64'h0593863e_4685fe04,
        64'h2783fef4_202337c1,
        64'h010007b7_4ee79f23,
        64'h47451ffe_b797998f,
        64'hf0effc84_350385be,
        64'hfc043603_2781fe64,
        64'h5783ffcf_f0ef853e,
        64'h4591863a_fe445703,
        64'h43dcfc84_3783fef4,
        64'h12238ff9_17fd6785,
        64'hfe445703_fef41223,
        64'h04000793_fef41323,
        64'h4785fce7_dee303f0,
        64'h07930007_871bfe84,
        64'h2783fef4_24232785,
        64'hfe842783_00078023,
        64'h97bafc04_3703fe84,
        64'h2783a235_478556e7,
        64'haa234705_1ffeb797,
        64'hd4dfc0ef_4f450513,
        64'h00001517_4ec58593,
        64'h00001597_1a000613,
        64'ha081fe04_24235807,
        64'had231ffe_b797a285,
        64'h47855ae7_a4234705,
        64'h1ffeb797_d81fc0ef,
        64'h52850513_00001517,
        64'h52058593_00001597,
        64'h19f00613_a02502f7,
        64'h1d631117_87931111,
        64'h17b7873e_53dcfc84,
        64'h37835c07_af231ffe,
        64'hb797c385_fc843783,
        64'hfcb43023_fca43423,
        64'h0080f822_fc067139,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aa851f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783911f,
        64'hf0ef853e_03e00593,
        64'h863a9341_1742fe84,
        64'h270343dc_fd843783,
        64'hfef42423_8fd9fe84,
        64'h278357f8_fd843783,
        64'hfef42423_8ff917e1,
        64'h67c1fe84_2703fef4,
        64'h242387aa_915ff0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_04f71963,
        64'h4791873e_57fcfd84,
        64'h37839edf_f0ef853e,
        64'h02800593_863a0ff7,
        64'h7713fe84_270343dc,
        64'hfd843783_fef42423,
        64'h0027e793_fe842783,
        64'ha039fef4_24230207,
        64'he793fe84_278300f7,
        64'h1963478d_873e0377,
        64'hc783fd84_3783fef4,
        64'h242387aa_9fdff0ef,
        64'h853e0280_059343dc,
        64'hfd843783_8c2fd0ef,
        64'h3e800513_9cfff0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe842783,
        64'ha8f5fef4_26234785,
        64'h9f3ff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe84,
        64'h2703fef4_242387aa,
        64'h9e1ff0ef_853e0300,
        64'h059343dc_fd843783,
        64'haa35fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa9d7f,
        64'he0effd84_35036000,
        64'h0593863e_4681fe44,
        64'h2783fef4_22231007,
        64'h879b03b7_07b7a039,
        64'hfef42223_5007879b,
        64'h03b707b7_00f71963,
        64'h4791873e_57fcfd84,
        64'h3783a02d_fef42223,
        64'h2007879b_03b707b7,
        64'ha825fef4_22236007,
        64'h879b03b7_07b700f7,
        64'h19634791_873e57fc,
        64'hfd843783_02f71763,
        64'h478d873e_0377c783,
        64'hfd843783_02e78ba3,
        64'h4709fd84_3783a031,
        64'h02e78ba3_470dfd84,
        64'h378300f7_186347a1,
        64'h873e4bdc_fd843783,
        64'h00f71f63_4795873e,
        64'h0347c783_fd843783,
        64'h02f71763_4789873e,
        64'h0367c783_fd843783,
        64'ha431fef4_26234785,
        64'h12078c63_2781fec4,
        64'h2783fef4_262387aa,
        64'haa9fe0ef_fd843503,
        64'h60078593_67a1863e,
        64'h4681fe44_2783fef4,
        64'h22230377_c783fd84,
        64'h378302e7_8ba34709,
        64'hfd843783_ac81fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaaebf_e0effd84,
        64'h35037007_8593678d,
        64'h863e4681_4bbcfd84,
        64'h378306f7_1b634785,
        64'h873e0347_c783fd84,
        64'h3783a479_fe042623,
        64'h00e7e563_478d873e,
        64'h4bdcfd84_3783a45d,
        64'h47858ae7_a8234705,
        64'h1ffec797_888fd0ef,
        64'h83050513_00002517,
        64'h82858593_00002597,
        64'h11300613_a02504f7,
        64'h10634789_873e0367,
        64'hc783fd84_37838e07,
        64'ha1231ffe_c797a4dd,
        64'h47858ee7_a8234705,
        64'h1ffec797_8c8fd0ef,
        64'h87050513_00002517,
        64'h86858593_00002597,
        64'h11200613_a02504f7,
        64'h13631117_87931111,
        64'h17b7873e_53dcfd84,
        64'h37839207_a3231ffe,
        64'hc797c385_fd843783,
        64'hfca43c23_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aab95f,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfd84,
        64'h3783c55f_f0ef853e,
        64'h03000593_460943dc,
        64'hfd843783_dfc52781,
        64'h8b89fe04_2783a83d,
        64'hfef42623_4785c79f,
        64'hf0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c3852781,
        64'h8ff967a1_fe042703,
        64'hfef42023_87aac67f,
        64'hf0ef853e_03000593,
        64'h43dcfd84_3783a8bd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_c5dfe0ef,
        64'hfd843503_30078593,
        64'h67ad4601_86be2781,
        64'hfe645783_9ee79f23,
        64'h47451ffe_c797e98f,
        64'hf0effd84_350385be,
        64'hfd043603_2781fe64,
        64'h5783cfdf_f0ef853e,
        64'h4591863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12238ff9_17fd6785,
        64'hfe445703_fef41223,
        64'h47a1fef4_13234785,
        64'ha8e5fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aacd7f,
        64'he0effd84_35037007,
        64'h8593678d_863e4681,
        64'h4bbcfd84_3783fce7,
        64'hdfe3479d_0007871b,
        64'hfe842783_fef42423,
        64'h2785fe84_27830007,
        64'h802397ba_fd043703,
        64'hfe842783_aa814785,
        64'ha8e7af23_47051ffe,
        64'hc797a76f_d0efa1e5,
        64'h05130000_2517a165,
        64'h85930000_25970ba0,
        64'h0613a081_fe042423,
        64'hac07a223_1ffec797,
        64'ha2514785_ace7a923,
        64'h47051ffe_c797aaaf,
        64'hd0efa525_05130000,
        64'h2517a4a5_85930000,
        64'h25970b90_0613a025,
        64'h02f71d63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_b007a423,
        64'h1ffec797_c385fd84,
        64'h3783fcb4_3823fca4,
        64'h3c231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_e1fff0ef,
        64'h85364591_863e93c1,
        64'h17c28ff9_17fd6785,
        64'hfd645703_43d4fd84,
        64'h3783fef4_26232781,
        64'h87aad99f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783a081,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_e05fe0ef,
        64'hfd843503_6585863e,
        64'h46812781_fd645783,
        64'ha0adfef4_26234785,
        64'ha89d4785_bae7a523,
        64'h47051ffe_c797b82f,
        64'hd0efb2a5_05130000,
        64'h2517b225_85930000,
        64'h259707f0_0613a025,
        64'hcb8d2781_3037f793,
        64'hfe842783_fef42423,
        64'h87aae19f_f0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'hbe07aa23_1ffec797,
        64'ha0f94785_c0e7a123,
        64'h47051ffe_c797bdaf,
        64'hd0efb825_05130000,
        64'h2517b7a5_85930000,
        64'h259707e0_0613a025,
        64'h04f71f63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_c207ac23,
        64'h1ffec797_c385fd84,
        64'h3783fcf4_1b2387ae,
        64'hfca43c23_1800f022,
        64'hf4067179_80826105,
        64'h644260e2_0001eb7f,
        64'hf0ef853e_85bafea4,
        64'h47039381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef40523,
        64'h87bafef4_05a387b6,
        64'hfef42623_873286ae,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e2853e_87aaea9f,
        64'hf0ef853e_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h05a387ba_fef42623,
        64'h872e87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_0001f63f,
        64'hf0ef853e_85bafe84,
        64'h57039381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef41423,
        64'h87bafef4_05a387b6,
        64'hfef42623_873286ae,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e2853e_87aaf47f,
        64'hf0ef853e_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h05a387ba_fef42623,
        64'h872e87aa_1000e822,
        64'hec061101_80826145,
        64'h74220001_00e79023,
        64'hfd645703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf41b23_87aefca4,
        64'h3c231800_f4227179,
        64'h80826145_74220001,
        64'h00e78023_fd744703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf40ba3,
        64'h87aefca4_3c231800,
        64'hf4227179_80826105,
        64'h6462853e_2781439c,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61056462_853e93c1,
        64'h17c20007_d783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826105,
        64'h6462853e_0ff7f793,
        64'h0007c783_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61616406,
        64'h60a6853e_fec42783,
        64'hfe042623_d3f8fb84,
        64'h37830007_871b0097,
        64'hd79bfd84_2783fcf4,
        64'h2c2302f7_07bbfe04,
        64'h2783fd84_2703fcf4,
        64'h2c2302f7_07bbfdc4,
        64'h27032781_2785fd84,
        64'h2783fcf4_2c238fd9,
        64'hfd842783_0007871b,
        64'h8ff9c007_87936785,
        64'h873e2781_00a7979b,
        64'hfd042783_fcf42c23,
        64'h0167d79b_fcc42783,
        64'hfcf42e23_278100f7,
        64'h17bb4705_27812789,
        64'h27818b9d_27810077,
        64'hd79bfcc4_2783fef4,
        64'h20232781_00f717bb,
        64'h47052781_8bbd2781,
        64'h0087d79b_fd042783,
        64'h02e78aa3_fb843783,
        64'h0ff7f713_8bbd0ff7,
        64'hf7932781_0127d79b,
        64'hfd442783_fcf42a23,
        64'h278187aa_9bdfd0ef,
        64'h853e9381_17822781,
        64'h27f143dc_fb843783,
        64'hfcf42823_278187aa,
        64'h9d9fd0ef_853e9381,
        64'h17822781_27e143dc,
        64'hfb843783_fcf42623,
        64'h278187aa_9f5fd0ef,
        64'h853e9381_17822781,
        64'h27d143dc_fb843783,
        64'hfcf42423_278187aa,
        64'ha11fd0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_a23dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa9d2f_f0effb84,
        64'h35039007_85936785,
        64'h863e4681_4bbcfb84,
        64'h3783aab1_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'ha00ff0ef_fb843503,
        64'h30000593_863e4681,
        64'h4bbcfb84_3783cbb8,
        64'h12340737_fb843783,
        64'hc7f8fb84_37830007,
        64'h871b87aa_b31fd0ef,
        64'h853e45f1_43dcfb84,
        64'h3783c7b8_fb843783,
        64'h0007871b_87aab4bf,
        64'hd0ef853e_45e143dc,
        64'hfb843783_c3f8fb84,
        64'h37830007_871b87aa,
        64'hb65fd0ef_853e45d1,
        64'h43dcfb84_3783c3b8,
        64'hfb843783_0007871b,
        64'h87aab7ff_d0ef853e,
        64'h45c143dc_fb843783,
        64'haaedfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaa9ef,
        64'hf0effb84_35032000,
        64'h05934601_4681db98,
        64'h4705fb84_3783c789,
        64'h27818ff9_400007b7,
        64'hfe842703_fa07dde3,
        64'hfe842783_fef42423,
        64'h87aab3bf_d0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783aca1,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_afcff0ef,
        64'hfb843503_10000593,
        64'h40ff8637_4681a091,
        64'hfe042423_a459fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aab2af_f0effb84,
        64'h35034581_46014681,
        64'ha46dfef4_26234785,
        64'he7892781_8ff967c1,
        64'hfe442703_fef42223,
        64'h87aabbbf_d0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fb843783,
        64'hcb8d47dc_fb843783,
        64'h02f70e63_400007b7,
        64'h873e2781_8ff9c000,
        64'h07b7873e_579cfb84,
        64'h3783a601_478510e7,
        64'haa234705_1ffec797,
        64'h8edfd0ef_07450513,
        64'h00002517_07458593,
        64'h00002597_67100613,
        64'ha02504f7_13634789,
        64'h873e0367_c783fb84,
        64'h37831407_a3231ffe,
        64'hc797a681_478514e7,
        64'haa234705_1ffec797,
        64'h92dfd0ef_0b450513,
        64'h00002517_0b458593,
        64'h00002597_67000613,
        64'ha02504f7_13631117,
        64'h87931111_17b7873e,
        64'h53dcfb84_37831807,
        64'ha5231ffe_c797c385,
        64'hfb843783_faa43c23,
        64'h0880e0a2_e486715d,
        64'h80826121_744270e2,
        64'h0001d05f_d0ef853a,
        64'h85be2781_08078793,
        64'hfd843783_93010207,
        64'h97132781_0587879b,
        64'h43dcfd84_378300e7,
        64'h912397b6_078e07c1,
        64'h93810206_1793fd84,
        64'h36839341_03079713,
        64'h02f707bb_0006861b,
        64'h36fdfec4_268393c1,
        64'h17c2fe44_27839341,
        64'h03079713_fd442783,
        64'h00e79023_02300713,
        64'h97ba078e_07c19381,
        64'h1782fd84_37032781,
        64'h37fdfec4_2783c3d8,
        64'h97b6078e_07c19381,
        64'h02061793_fd843683,
        64'h0007871b_9fb90006,
        64'h861b36fd_fec42683,
        64'h27810107_979bfe84,
        64'h27830007_871bfc84,
        64'h3783f8e7_ebe32781,
        64'hfe842783_0007871b,
        64'h37fdfec4_2783fef4,
        64'h24232785_fe842783,
        64'h00079123_97ba078e,
        64'h07c1fe84_6783fd84,
        64'h370300e7_90230210,
        64'h071397ba_078e07c1,
        64'hfe846783_fd843703,
        64'hc3d897b6_078e07c1,
        64'hfe846783_fd843683,
        64'h0007871b_9fb92781,
        64'h0107979b_fe842783,
        64'h0007871b_fc843783,
        64'ha8b1fe04_2423fef4,
        64'h26232785_fec42783,
        64'hc7912781_8ff917fd,
        64'h67c1873e_278102f7,
        64'h07bbfe44_2783fd44,
        64'h2703fef4_26230107,
        64'hd79b2781_02f707bb,
        64'hfe442783_fd442703,
        64'ha835fef4_26234785,
        64'h00f77663_67c1873e,
        64'h278102f7_07bbfe44,
        64'h2783fd44_2703fef4,
        64'h22238ff9_17fd6785,
        64'hfe442703_fef42223,
        64'h87aaebff_d0ef853e,
        64'h459143dc_fd843783,
        64'hfe042223_fe042423,
        64'hfe042623_fcf42a23,
        64'hfcc43423_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_61457402,
        64'h70a2853e_fec42783,
        64'h0001a011_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'he10ff0ef_fd843503,
        64'h70000593_863e4681,
        64'h4bbcfd84_3783fe04,
        64'h2623fca4_3c231800,
        64'hf022f406_71798082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hf87fd0ef_853e0300,
        64'h05934609_43dcfd84,
        64'h3783dfc5_27818b89,
        64'hfe442783_a00dfef4,
        64'h26234785_fabfd0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_f99fd0ef,
        64'h853e0300_059343dc,
        64'hfd843783_a08dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaebaf_f0effd84,
        64'h35039007_85936789,
        64'h863e86ba_fd442783,
        64'hfd042703_46e79023,
        64'h02700713_1ffec797,
        64'ha879fef4_26234785,
        64'hc3b92781_fec42783,
        64'hfef42623_87aaef6f,
        64'hf0effd84_35038007,
        64'h85936789_863e86ba,
        64'hfd442783_fd042703,
        64'h48e79d23_470d1ffe,
        64'hc79702f7_1f634785,
        64'h0007871b_fd042783,
        64'h142000ef_fd843503,
        64'h85befc84_3603fd04,
        64'h2783a8e5_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h081000ef_fd843503,
        64'h20000593_02f70363,
        64'h20000793_873e2781,
        64'h87aafd3f_d0ef853e,
        64'h93811782_27812791,
        64'h43dcfd84_3783aa35,
        64'hfef42623_4785e789,
        64'h27818ff9_67c1fe84,
        64'h2703fef4_242387aa,
        64'h800fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783cb8d,
        64'h47dcfd84_378302f7,
        64'h0e634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_fd843783,
        64'h00f71f63_4789873e,
        64'h0367c783_fd843783,
        64'hfcf42823_87bafcf4,
        64'h2a23fcd4_34238732,
        64'h87aefca4_3c230080,
        64'hf822fc06_71398082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'h880fe0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_96afe0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe442783,
        64'ha83dfef4_26234785,
        64'h98efe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe44,
        64'h2703fef4_222387aa,
        64'h97cfe0ef_853e0300,
        64'h059343dc_fd843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa89ff,
        64'hf0effd84_35032007,
        64'h85936785_863e86ba,
        64'hfd442783_fd042703,
        64'h64e79223_03700713,
        64'h1ffec797_a86dfef4,
        64'h26234785_c3b92781,
        64'hfec42783_fef42623,
        64'h87aa8dbf_f0effd84,
        64'h35031007_85936785,
        64'h863e86ba_fd442783,
        64'hfd042703_66e79f23,
        64'h474d1ffe_c79702f7,
        64'h1f634785_0007871b,
        64'hfd042783_326000ef,
        64'hfd843503_85befc84,
        64'h3603fd04_2783aa11,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_265000ef,
        64'hfd843503_20000593,
        64'h02f70363_20000793,
        64'h873e2781_87aa9b6f,
        64'he0ef853e_93811782,
        64'h27812791_43dcfd84,
        64'h3783aaa1_fef42623,
        64'h4785e789_27818ff9,
        64'h67c1fe84_2703fef4,
        64'h242387aa_9e4fe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783cb8d_47dcfd84,
        64'h378302f7_0e634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfd843783_00f71f63,
        64'h4789873e_0367c783,
        64'hfd843783_fcf42823,
        64'h87bafcf4_2a23fcd4,
        64'h34238732_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_61457422,
        64'h853efec4_27830001,
        64'ha0110001_a0210001,
        64'ha031fef4_26238fd9,
        64'hfd442783_fec42703,
        64'ha831fef4_262301a7,
        64'he793fec4_2783a02d,
        64'hfef42623_03a7e793,
        64'hfec42783_a825fef4,
        64'h262301a7_e793fec4,
        64'h2783a099_fef42623,
        64'h0027e793_fec42783,
        64'ha891fef4_262303a7,
        64'he793fec4_2783a08d,
        64'hfef42623_03a7e793,
        64'hfec42783_a885fef4,
        64'h262301a7_e793fec4,
        64'h2783a8bd_fef42623,
        64'h0097e793_fec42783,
        64'ha071fef4_262303a7,
        64'he793fec4_2783a869,
        64'hfef42623_01a7e793,
        64'hfec42783_00f71963,
        64'h4785873e_0347c783,
        64'hfd843783_a865fef4,
        64'h262301a7_e793fec4,
        64'h2783a0d9_fef42623,
        64'h01a7e793_fec42783,
        64'ha8d1fef4_262301b7,
        64'he793fec4_2783a0cd,
        64'hfef42623_03a7e793,
        64'hfec42783_00f71963,
        64'h4785873e_0347c783,
        64'hfd843783_a201fef4,
        64'h262301b7_e793fec4,
        64'h2783a239_fef42623,
        64'h01b7e793_fec42783,
        64'haa31fef4_26230097,
        64'he793fec4_2783a22d,
        64'hfef42623_0027e793,
        64'hfec42783_aa390ef7,
        64'h05639007_879367ad,
        64'h0007871b_10e68a63,
        64'h30070713_672d0007,
        64'h869b10e6_8a63a007,
        64'h0713672d_0007869b,
        64'ha2a916f7_0363a007,
        64'h87936791_0007871b,
        64'h0ee68d63_d0070713,
        64'h67250007_869b0ae6,
        64'h89636007_07136721,
        64'h0007869b_02d76863,
        64'h70070713_67250007,
        64'h869b14e6_80637007,
        64'h07136725_0007869b,
        64'haa4914f7_08638007,
        64'h87936789_0007871b,
        64'h18e68b63_40070713,
        64'h670d0007_869b16e6,
        64'h86639007_07136709,
        64'h0007869b_aa7d16f7,
        64'h07632007_87936785,
        64'h0007871b_16e68e63,
        64'h50070713_67050007,
        64'h869b18e6_85633007,
        64'h07136705_0007869b,
        64'h02d76863_70070713,
        64'h67050007_869b1ae6,
        64'h8a637007_07136705,
        64'h0007869b_06d76c63,
        64'h70070713_670d0007,
        64'h869b20e6_84637007,
        64'h0713670d_0007869b,
        64'ha40d1cf7_0263b007,
        64'h87936785_0007871b,
        64'h1ce68963_67050007,
        64'h869b1ce6_8e63c007,
        64'h07136705_0007869b,
        64'ha4a91af7_02637000,
        64'h07930007_871b1ee6,
        64'h85639007_07136705,
        64'h0007869b_1c070663,
        64'h27018007_871b02d7,
        64'h6563a007_07136705,
        64'h0007869b_20e68f63,
        64'ha0070713_67050007,
        64'h869ba471_18f70863,
        64'h30000793_0007871b,
        64'h1ae68563_50000713,
        64'h0007869b_2ae68e63,
        64'h40000713_0007869b,
        64'hac4d18f7_0d631000,
        64'h07930007_871b2c07,
        64'h09630007_871b00d7,
        64'h6d632000_07130007,
        64'h869b1ce6_84632000,
        64'h07130007_869b04d7,
        64'h6c636000_07130007,
        64'h869b20e6_85636000,
        64'h07130007_869b0cd7,
        64'h6d631007_07136705,
        64'h0007869b_2ae68a63,
        64'h10070713_67050007,
        64'h869bfd44_2783fef4,
        64'h2623fd44_2783fcf4,
        64'h2a2387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'he86fe0ef_853e0300,
        64'h05934605_43dcfd84,
        64'h3783d3a9_27818b85,
        64'hfe042783_a00dea4f,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_fef42623,
        64'h4789e781_27819bf9,
        64'hfec42783_fef42623,
        64'h87aae96f_e0ef853e,
        64'h03200593_43dcfd84,
        64'h3783c3a1_27818ff9,
        64'h67a1fe04_2703a899,
        64'heeefe0ef_853e0300,
        64'h05930200_061343dc,
        64'hfd843783_cf812781,
        64'h0207f793_278187aa,
        64'hed4fe0ef_853e0300,
        64'h059343dc_fd843783,
        64'h02f71b63_30078793,
        64'h67850007_871bfd44,
        64'h278300f7_0b635007,
        64'h87936785_0007871b,
        64'hfd442783_fef42023,
        64'h87aaf0ef_e0ef853e,
        64'h03000593_43dcfd84,
        64'h3783ef4f_e0ef853a,
        64'h85be2781_8fd52781,
        64'hbb07d783_1ffed797,
        64'h0007869b_0107979b,
        64'hfe442783_93010207,
        64'h97132781_27b143dc,
        64'hfd843783_a229fef4,
        64'h26234785_c7892781,
        64'h0207f793_fe442783,
        64'hcb992781_8b89fe84,
        64'h2783fef4_242387aa,
        64'hed8fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_378302f7,
        64'h0f633007_87936785,
        64'h0007871b_fd442783,
        64'h04f70863_50078793,
        64'h67850007_871bfd44,
        64'h2783fef4_22238ff9,
        64'h17fd6791_fe442703,
        64'hfef42223_87aa18c0,
        64'h00effd84_350385be,
        64'hfd442783_80bfe0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783821f_e0ef853a,
        64'h03000593_fff78613,
        64'h67c143d8_fd843783,
        64'hfd2fe0ef_853e85ba,
        64'hfd042703_93811782,
        64'h278127a1_43dcfd84,
        64'h37838d1f_e0ef853e,
        64'h02e00593_463943dc,
        64'hfd843783_863fe0ef,
        64'h853e4599_863a9341,
        64'h1742fcc4_270343dc,
        64'hfd843783_aaedfef4,
        64'h26234785_a4194785,
        64'hcce7a723_47051ffe,
        64'hd797ca6f_e0efc2e5,
        64'h05130000_3517c2e5,
        64'h85930000_359744c0,
        64'h0613a025_cb8d2781,
        64'h8b85fe84_2783fef4,
        64'h242387aa_fe4fe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783d007_ab231ffe,
        64'hd797acb1_4785d2e7,
        64'ha2234705_1ffed797,
        64'hcfcfe0ef_c8450513,
        64'h00003517_c8458593,
        64'h00003597_44b00613,
        64'ha02504f7_1e631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783d407,
        64'had231ffe_d797c385,
        64'hfd843783_fcf42623,
        64'h87bafcf4_282387b2,
        64'hfcf42a23_873687ae,
        64'hfca43c23_0080f822,
        64'hfc067139_80826145,
        64'h740270a2_853efec4,
        64'h27830001_fcf719e3,
        64'h01f007b7_873e2781,
        64'h8ff901f0_07b7fe84,
        64'h2703fef4_242387aa,
        64'h899fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783a839,
        64'hfef42423_87aa8b7f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_fcafe0ef,
        64'h3e800513_9abfe0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0047e793,
        64'h93c117c2_fe442783,
        64'h43d8fd84_3783fef4,
        64'h222387aa_999fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_d3ed2781,
        64'h8b89fe44_2783fef4,
        64'h222387aa_9b9fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a821fef4,
        64'h222387aa_9d1fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a1bfe0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0017e793,
        64'h93c117c2_fe442783,
        64'h43d8fd84_3783fef4,
        64'h222387aa_a09fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a211fef4,
        64'h26234785_e7892781,
        64'h8ba12781_fe245783,
        64'hfef41123_87aaa33f,
        64'he0ef853e_03e00593,
        64'h43dcfd84_37838a5f,
        64'he0ef3887_85136785,
        64'ha87fe0ef_853e03e0,
        64'h0593863a_fe245703,
        64'h43dcfd84_3783fef4,
        64'h11230087_e793fe24,
        64'h5783fef4_112387aa,
        64'ha75fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'habffe0ef_853e02c0,
        64'h0593863a_fe245703,
        64'h43dcfd84_3783fef4,
        64'h11239be9_fe245783,
        64'hfef41123_87aaaabf,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783ffe1,
        64'h27818ff9_01f007b7,
        64'hfe842703_fef42423,
        64'h87aaa33f_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'ha839fef4_242387aa,
        64'ha51fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783fef4,
        64'h26234785_c7812781,
        64'hfec42783_fef42623,
        64'h87aa2120_00effd84,
        64'h3503b007_85936785,
        64'h46014681_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623f3e5_27818b89,
        64'h2781feb4_4783fef4,
        64'h05a387aa_bd9fe0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_a821fef4,
        64'h05a387aa_bf1fe0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_c3bfe0ef,
        64'h853e02f0_05934609,
        64'h43dcfd84_3783bcdf,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_be3fe0ef,
        64'h853a0300_0593fff7,
        64'h861367c1_43d8fd84,
        64'h378302e7_8a234709,
        64'hfd843783_a03102e7,
        64'h8a234705_fd843783,
        64'hc7992781_fec42783,
        64'hfef42623_87aa2de0,
        64'h00effd84_35031000,
        64'h059340ff_86374681,
        64'ha855fef4_26234785,
        64'ha0c14785_08e7a123,
        64'h47051ffe_d79785bf,
        64'he0effe25_05130000,
        64'h3517fe25_85930000,
        64'h35973ac0_0613a025,
        64'hcb8d2781_fec42783,
        64'hfef42623_87aa32e0,
        64'h00effd84_35034581,
        64'h46014681_aa3fe0ef,
        64'h71078513_67890c07,
        64'ha5231ffe_d797aa19,
        64'h47850ce7_ac234705,
        64'h1ffed797_8b1fe0ef,
        64'h03850513_00003517,
        64'h03858593_00003597,
        64'h3ab00613_a02504f7,
        64'h1e631117_87931111,
        64'h17b7873e_53dcfd84,
        64'h37831007_a7231ffe,
        64'hd797c385_fd843783,
        64'hfca43c23_1800f022,
        64'hf4067179_8082614d,
        64'h64ea740a_70aa853e,
        64'hfdc42783_0001a011,
        64'h0001a021_0001a031,
        64'hfcf42e23_4785cb89,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_504010ef,
        64'hf5843503_20000593,
        64'h02f71763_4785873e,
        64'h0347c783_f5843783,
        64'h00f71a63_4791873e,
        64'h57fcf584_37830001,
        64'ha0b9fcf4_2e234785,
        64'hc7912781_fdc42783,
        64'hfcf42e23_87aa79e0,
        64'h20eff584_350385be,
        64'hfd442783_fcf42a23,
        64'h1007879b_03a207b7,
        64'heb950a27_c783fb67,
        64'h87931ffe_d797a071,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_09d010ef,
        64'hf5843503_02f71163,
        64'h4791873e_57fcf584,
        64'h3783a865_fcf42e23,
        64'h478500f7_06634785,
        64'h873e0b97_c783ffe7,
        64'h87931ffe_d79704f7,
        64'h16634791_873e57fc,
        64'hf5843783_00f70963,
        64'h4795873e_57fcf584,
        64'h3783a8c5_fcf42e23,
        64'h478500f7_06634789,
        64'h873e0b97_c7830367,
        64'h87931ffe_d79702f7,
        64'h1063479d_873e57fc,
        64'hf5843783_aa29fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa6ac0_20eff584,
        64'h350306a5_85931ffe,
        64'hd597a281_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h657010ef_f5843503,
        64'h0cf70b63_4799873e,
        64'h57fcf584_3783d7f8,
        64'h4719f584_3783a029,
        64'hd7f84715_f5843783,
        64'h00e7f763_4785873e,
        64'h0377c783_f5843783,
        64'hcf912781_8b892781,
        64'h0c47c783_0cc78793,
        64'h1ffed797_a825d7f8,
        64'h4711f584_378300e7,
        64'hf7634785_873e0377,
        64'hc783f584_3783cf91,
        64'h27818bb1_27810c47,
        64'hc7830fa7_87931ffe,
        64'hd797a09d_d7f8471d,
        64'hf5843783_00e7f763,
        64'h4785873e_0377c783,
        64'hf5843783_cf912781,
        64'h0307f793_27810c47,
        64'hc78312a7_87931ffe,
        64'hd797d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0d47c783_14478793,
        64'h1ffed797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0087979b_27810d57,
        64'hc78316a7_87931ffe,
        64'hd79753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810107,
        64'h979b2781_0d67c783,
        64'h19078793_1ffed797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h0187979b_27810d77,
        64'hc7831b27_87931ffe,
        64'hd797a461_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h01b020ef_f5843503,
        64'h1d858593_1ffed597,
        64'ha47dfcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa2bf0,
        64'h10eff584_350328f7,
        64'h12634795_873e0347,
        64'hc783f584_3783acf1,
        64'hfcf42e23_478528f7,
        64'h0d634785_873e0b97,
        64'hc7832227_87931ffe,
        64'hd797ace5_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h08b020ef_f5843503,
        64'h24858593_1ffed597,
        64'hae39fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa0340,
        64'h20eff584_3503d7f8,
        64'h4715f584_37832ee7,
        64'hfd634785_873e0377,
        64'hc783f584_37833007,
        64'h85632781_8b892781,
        64'h0c47c783_29478793,
        64'h1ffed797_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810d47_c7832ae7,
        64'h87931ffe_d79753f8,
        64'hf5843783_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810087_979b2781,
        64'h0d57c783_2d478793,
        64'h1ffed797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0107979b_27810d67,
        64'hc7832fa7_87931ffe,
        64'hd79753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b0187_979b2781,
        64'h0d77c783_31c78793,
        64'h1ffed797_aecdfcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa1850_20eff584,
        64'h35033425_85931ffe,
        64'hd597a921_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h429010ef_f5843503,
        64'h14f71f63_4785873e,
        64'h0367c783_f5843783,
        64'h16e7f763_478d873e,
        64'h0357c783_f5843783,
        64'h16f71f63_4789873e,
        64'h0347c783_f5843783,
        64'ha19dfcf4_2e234785,
        64'h42078363_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h17e020ef_f5843503,
        64'hd7f84715_f5843783,
        64'h44e7f363_4785873e,
        64'h0377c783_f5843783,
        64'h44078b63_27818b89,
        64'h2781f9d4_47834607,
        64'h82630004_c78302e7,
        64'h8e234705_f5843783,
        64'hfd7fe0ef_3e800513,
        64'h9b6ff0ef_853a02c0,
        64'h0593863e_93c117c2,
        64'h0047e793_fda45783,
        64'h43d8f584_3783fcf4,
        64'h1d2387aa_9a0ff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_d3e52781,
        64'h8b892781_fda45783,
        64'hfcf41d23_87aa9c2f,
        64'hf0ef853e_02c00593,
        64'h43dcf584_3783a821,
        64'hfcf41d23_87aa9daf,
        64'hf0ef853e_02c00593,
        64'h43dcf584_3783a24f,
        64'hf0ef853a_02c00593,
        64'h863e93c1_17c20017,
        64'he793fda4_578343d8,
        64'hf5843783_fcf41d23,
        64'h87aaa0ef_f0ef853e,
        64'h02c00593_43dcf584,
        64'h3783a3a5_fcf42e23,
        64'h4785e789_27818ba1,
        64'h2781fd24_5783fcf4,
        64'h192387aa_a38ff0ef,
        64'h853e03e0_059343dc,
        64'hf5843783_8aaff0ef,
        64'h38878513_6785a8cf,
        64'hf0ef853e_03e00593,
        64'h863afd24_570343dc,
        64'hf5843783_fcf41923,
        64'h0087e793_fd245783,
        64'hfcf41923_87aaa7af,
        64'hf0ef853e_03e00593,
        64'h43dcf584_3783ac4f,
        64'hf0ef853e_02c00593,
        64'h863afd24_570343dc,
        64'hf5843783_fcf41923,
        64'h9be9fd24_5783fcf4,
        64'h192387aa_ab0ff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_14079d63,
        64'h03c7c783_f5843783,
        64'h16f71363_47a1873e,
        64'h4bdcf584_378316e7,
        64'hfa63478d_873ef9d4,
        64'h47831807_d0634187,
        64'hd79b0187_979b0024,
        64'hc7836207_9e632781,
        64'hfdc42783_fcf42e23,
        64'h87aa18e0_20eff584,
        64'h350385be_f9040793,
        64'hadb9fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa66f0,
        64'h10eff584_3503c385,
        64'h27818b91_27810014,
        64'hc783a561_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h4b3010ef_f5843503,
        64'h85a6a565_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h34d020ef_f5843503,
        64'h26f71263_4785873e,
        64'h0347c783_f5843783,
        64'hadd9fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa46c0,
        64'h10eff584_3503add5,
        64'hfcf42e23_4785adf5,
        64'hfcf42e23_4785cb89,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_06f020ef,
        64'hf5843503_85be5f9c,
        64'hf5843783_df98a807,
        64'h071b018c_c737f584,
        64'h3783af05_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h6dc010ef_f5843503,
        64'h04f71b63_4795873e,
        64'h0347c783_f5843783,
        64'h00f70a63_4789873e,
        64'h0347c783_f5843783,
        64'ha7bdfcf4_2e234785,
        64'hc3d12781_fdc42783,
        64'hfcf42e23_87aa0e10,
        64'h20eff584_350385be,
        64'h5f9cf584_3783df98,
        64'h8407071b_017d8737,
        64'hf5843783_a801df98,
        64'hac07071b_0121f737,
        64'hf5843783_00f71a63,
        64'h4789873e_0367c783,
        64'hf5843783_7c40006f,
        64'hfcf42e23_4785c791,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_915ff0ef,
        64'hf5843503_06f71c63,
        64'h4785873e_0347c783,
        64'hf5843783_7f40006f,
        64'hfcf42e23_478500f7,
        64'h07634795_873e0347,
        64'hc783f584_378300f7,
        64'h0f634789_873e0347,
        64'hc783f584_378302f7,
        64'h07634785_873e0347,
        64'hc783f584_378302f7,
        64'h02e34785_0007871b,
        64'hfdc42783_fcf42e23,
        64'h87aa0530_00eff584,
        64'h3503a839_02e78a23,
        64'h4715f584_378300f7,
        64'h18634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_f5843783,
        64'h0750006f_47859ae7,
        64'ha6234705_1ffee797,
        64'h984ff0ef_90c50513,
        64'h00004517_90c58593,
        64'h00004597_24000613,
        64'ha02d04f7_1a634789,
        64'h873e0367_c783f584,
        64'h3783df98_a807071b,
        64'h00062737_f5843783,
        64'h02078e23_f5843783,
        64'h02e78a23_4705f584,
        64'h378302e7_8ba34705,
        64'hf5843783_a007a423,
        64'h1ffee797_0e10006f,
        64'h4785a0e7_ac234705,
        64'h1ffee797_9f0ff0ef,
        64'h97850513_00004517,
        64'h97858593_00004597,
        64'h23f00613_a02d06f7,
        64'h19631117_87931111,
        64'h17b7873e_53dcf584,
        64'h3783a407_a7231ffe,
        64'he797c385_f5843783,
        64'hfc043423_fc043023,
        64'hfa043c23_fa043823,
        64'hfa043423_fa043023,
        64'hf8043c23_f8043823,
        64'h0004b023_00579493,
        64'h839507fd_f8078793,
        64'hfe040793_f4a43c23,
        64'h1900ed26_f122f506,
        64'h71718082_61616406,
        64'h60a6853e_fec42783,
        64'hfe042623_d3f8fb84,
        64'h37830007_871b00a7,
        64'h979b2781_27852781,
        64'h8ff917fd_004007b7,
        64'h873e2781_0087d79b,
        64'hfc442783_02f71663,
        64'h4785873e_27818b8d,
        64'h27810167_d79bfcc4,
        64'h2783a081_d3f8fb84,
        64'h37830007_871b0097,
        64'hd79bfd04_2783fcf4,
        64'h282302f7_07bbfd84,
        64'h2783fd04_2703fcf4,
        64'h282302f7_07bbfd44,
        64'h27032781_2785fd04,
        64'h2783fcf4_28238fd9,
        64'hfd042783_0007871b,
        64'h8ff9c007_87936785,
        64'h873e2781_00a7979b,
        64'hfc842783_fcf42823,
        64'h0167d79b_fc442783,
        64'hfcf42a23_278100f7,
        64'h17bb4705_27812789,
        64'h27818b9d_27810077,
        64'hd79bfc44_2783fcf4,
        64'h2c232781_00f717bb,
        64'h47052781_8bbd2781,
        64'h0087d79b_fc842783,
        64'he3c52781_8b8d2781,
        64'h0167d79b_fcc42783,
        64'hfcf42623_278187aa,
        64'he88ff0ef_853e9381,
        64'h17822781_27f143dc,
        64'hfb843783_fcf42423,
        64'h278187aa_ea4ff0ef,
        64'h853e9381_17822781,
        64'h27e143dc_fb843783,
        64'hfcf42223_278187aa,
        64'hec0ff0ef_853e9381,
        64'h17822781_27d143dc,
        64'hfb843783_fcf42023,
        64'h278187aa_edcff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'ha28dfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa69f0,
        64'h00effb84_35039007,
        64'h85936785_863e4681,
        64'h4bbcfb84_3783d7d5,
        64'h4bbcfb84_3783cbb8,
        64'hfb843783_0007871b,
        64'h8ff977c1_873e2781,
        64'h87aaf3af_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783a2c1,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_6fd000ef,
        64'hfb843503_30000593,
        64'h46014681_c7f8fb84,
        64'h37830007_871b87aa,
        64'h81dff0ef_853e45f1,
        64'h43dcfb84_3783c7b8,
        64'hfb843783_0007871b,
        64'h87aa837f_f0ef853e,
        64'h45e143dc_fb843783,
        64'hc3f8fb84_37830007,
        64'h871b87aa_851ff0ef,
        64'h853e45d1_43dcfb84,
        64'h3783c3b8_fb843783,
        64'h0007871b_87aa86bf,
        64'hf0ef853e_45c143dc,
        64'hfb843783_a4b9fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa78b0_00effb84,
        64'h35032000_05934601,
        64'h4681ac95_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h585000ef_fb843503,
        64'h02e78e23_4705fb84,
        64'h3783c78d_27818ff9,
        64'h010007b7_fe842703,
        64'hdb984705_fb843783,
        64'hc7892781_8ff94000,
        64'h07b7fe84_2703f407,
        64'hdde3fe84_2783fef4,
        64'h242387aa_85dff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'ha4cdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa01e0,
        64'h10effb84_35039007,
        64'h859367ad_863e4681,
        64'hfe442783_fef42223,
        64'h8fd90100_07b7fe44,
        64'h270300f7_196347a1,
        64'h873e4bdc_fb843783,
        64'h02f71063_4789873e,
        64'h0367c783_fb843783,
        64'hfef42223_40ff87b7,
        64'ha689fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa07e0,
        64'h10effb84_35037007,
        64'h8593678d_46014681,
        64'ha055fe04_242302e7,
        64'h8aa34709_fb843783,
        64'ha03102e7_8aa34705,
        64'hfb843783_00f70863,
        64'h1aa00793_0007871b,
        64'hfe842783_fef42423,
        64'h87aa92bf_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783f3e5,
        64'h27818b89_2781fe34,
        64'h4783fef4_01a387aa,
        64'ha6dff0ef_853e02f0,
        64'h059343dc_fb843783,
        64'ha821fef4_01a387aa,
        64'ha85ff0ef_853e02f0,
        64'h059343dc_fb843783,
        64'hacfff0ef_853e02f0,
        64'h05934609_43dcfb84,
        64'h378304f7_18634789,
        64'h0007871b_fec42783,
        64'ha129fef4_26234785,
        64'h00f70663_47890007,
        64'h871bfec4_2783cf81,
        64'h2781fec4_2783fef4,
        64'h262387aa_154010ef,
        64'hfb843503_80078593,
        64'h67851aa0_06134681,
        64'ha189fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa17e0,
        64'h10effb84_35034581,
        64'h46014681_a19dfef4,
        64'h26234785_e7892781,
        64'h8ff967c1_fdc42703,
        64'hfcf42e23_87aaa0ff,
        64'hf0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfb843783_cb8d47dc,
        64'hfb843783_02f70e63,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cfb84_3783a975,
        64'h4785f6e7_a4234705,
        64'h1ffee797_f40ff0ef,
        64'hec850513_00004517,
        64'hec858593_00004597,
        64'h16200613_a02504f7,
        64'h13634789_873e0367,
        64'hc783fb84_3783cbd8,
        64'h4711fb84_3783fa07,
        64'ha1231ffe_e797a311,
        64'h4785fae7_a8234705,
        64'h1ffee797_f88ff0ef,
        64'hf1050513_00004517,
        64'hf1058593_00004597,
        64'h16100613_a02504f7,
        64'h17631117_87931111,
        64'h17b7873e_53dcfb84,
        64'h3783fe07_a3231ffe,
        64'he797c385_fb843783,
        64'hfaa43c23_0880e0a2,
        64'he486715d_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623bcdf,
        64'hf0ef853e_45912000,
        64'h061343dc_fd843783,
        64'h02e79523_474d1ffe,
        64'he797be9f_f0ef853e,
        64'h03a00593_460143dc,
        64'hfd843783_bfbff0ef,
        64'h853e0380_05934601,
        64'h43dcfd84_3783c0df,
        64'hf0ef853a_03600593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c23ff0ef,
        64'h853a0340_0593eff7,
        64'h861367c1_43d8fd84,
        64'h3783cb9f_f0ef853e,
        64'h02800593_464143dc,
        64'hfd843783_ccbff0ef,
        64'h853a0290_0593863e,
        64'h0ff7f793_0017e793,
        64'hfeb44783_43d8fd84,
        64'h3783fe04_05a3a019,
        64'hfef405a3_47a9c789,
        64'h27818ff9_040007b7,
        64'h873e579c_fd843783,
        64'ha005fef4_05a347b1,
        64'hc7892781_8ff90200,
        64'h07b7873e_579cfd84,
        64'h3783a82d_fef405a3,
        64'h47b9c789_27818ff9,
        64'h010007b7_873e579c,
        64'hfd843783_a8d5fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa13c0_30effd84,
        64'h3503a807_85930006,
        64'h27b7b09f_f0ef0c80,
        64'h051300f7_16634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfd843783_02f71363,
        64'h4789873e_0367c783,
        64'hfd843783_d93ff0ef,
        64'h853e0290_0593463d,
        64'h43dcfd84_3783a811,
        64'hda7ff0ef_853e0290,
        64'h0593463d_43dcfd84,
        64'h378300f7_1c634789,
        64'h873e0367_c783fd84,
        64'h3783d798_fd843783,
        64'h0007871b_87aac7ff,
        64'hf0ef853e_93811782,
        64'h27810407_879b43dc,
        64'hfd843783_02e78b23,
        64'hfd843783_0ff7f713,
        64'h87aad3ff_f0ef853e,
        64'h0fe00593_43dcfd84,
        64'h3783f3e5_27818b85,
        64'h2781fea4_4783fef4,
        64'h052387aa_de1ff0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_a821fef4,
        64'h052387aa_df9ff0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_e43ff0ef,
        64'h853e02f0_05934605,
        64'h43dcfd84_3783bfdf,
        64'hf0ef3e80_0513e5df,
        64'hf0ef853e_02900593,
        64'h460143dc_fd843783,
        64'ha811e71f_f0ef853e,
        64'h02900593_464143dc,
        64'hfd843783_a4814785,
        64'h24e7a723_47051ffe,
        64'he797a27f_f0ef1ae5,
        64'h05130000_45171ae5,
        64'h85930000_45970b50,
        64'h0613a025_04f71063,
        64'h4789873e_27810ff7,
        64'hf7932781_87aae03f,
        64'hf0ef853e_0fe00593,
        64'h43dcfd84_37830607,
        64'hb823fd84_3783d7f8,
        64'h4719fd84_37830607,
        64'ha223fd84_378302e7,
        64'h8023fd84_37830207,
        64'hc703fd04_3783cfd8,
        64'hfd843783_4fd8fd04,
        64'h3783cf98_fd843783,
        64'h4f98fd04_3783cbd8,
        64'hfd843783_4bd8fd04,
        64'h3783cb98_fd843783,
        64'h4b98fd04_3783c7d8,
        64'hfd843783_47d8fd04,
        64'h3783d3d8_1117071b,
        64'h11111737_fd843783,
        64'hc798fd84_37834798,
        64'hfd043783_c3d8fcc4,
        64'h2703fd84_378300e7,
        64'h9023fd84_37830007,
        64'hd703fd04_37833207,
        64'ha5231ffe_e797a62d,
        64'h478532e7_ac234705,
        64'h1ffee797_b11ff0ef,
        64'h29850513_00004517,
        64'h29858593_00004597,
        64'h0b400613_a025c7fd,
        64'hfd043783_3607a023,
        64'h1ffee797_cb89fd84,
        64'h3783fcf4_262387b2,
        64'hfcb43823_fca43c23,
        64'h0080f822_fc067139,
        64'h80826105_644260e2,
        64'h0001e8df_f0ef853e,
        64'h85bafea4_47039381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef40523_87bafef4,
        64'h05a387b6_fef42623,
        64'h873286ae_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e2853e,
        64'h87aae7ff_f0ef853e,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_05a387ba,
        64'hfef42623_872e87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h0001f39f_f0ef853e,
        64'h85bafe84_57039381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef41423_87bafef4,
        64'h05a387b6_fef42623,
        64'h873286ae_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e2853e,
        64'h87aaf1df_f0ef853e,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_05a387ba,
        64'hfef42623_872e87aa,
        64'h1000e822_ec061101,
        64'h80826145_74220001,
        64'hc398fd44_2703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_2a2387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61457422,
        64'h000100e7_9023fd64,
        64'h5703fe84_3783fef4,
        64'h3423fd84_3783fcf4,
        64'h1b2387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61457422_000100e7,
        64'h8023fd74_4703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_0ba387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61056462,
        64'h853e2781_439cfe84,
        64'h3783fea4_34231000,
        64'hec221101_80826105,
        64'h6462853e_93c117c2,
        64'h0007d783_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61056462,
        64'h853e0ff7_f7930007,
        64'hc783fe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826145_7422853e,
        64'hfe843783_fae7f5e3,
        64'h47850007_871bfe44,
        64'h2783fef4_22232785,
        64'hfe442783_a829fef4,
        64'h342397ba_10470713,
        64'h00005717_078a97ba,
        64'h078e87ba_fe446703,
        64'h02f71063_27812701,
        64'hfde45703_0007d783,
        64'h97ba1366_8713078a,
        64'h97ba078e_87bafe44,
        64'h67030000_5697a0b9,
        64'hfe042223_fe043423,
        64'hfcf41f23_87aa1800,
        64'hf4227179_80826145,
        64'h740270a2_0001fef7,
        64'h68e3fe04_3783fe84,
        64'h3703fea4_3423fbff,
        64'hf0effef4_302397ba,
        64'hfe843783_873e078a,
        64'h97ba078a_87bafd84,
        64'h3703fea4_3423fdff,
        64'hf0effca4_3c231800,
        64'hf022f406_71798082,
        64'h01416422_853e639c,
        64'h17e10200_c7b70800,
        64'he4221141_80826109,
        64'h640660a6_853efec4,
        64'h2783fef4_262387aa,
        64'hb38ff0ef_c2650513,
        64'hfffff517_85be567d,
        64'hfb843683_fd040793,
        64'hfe043703_fcf43c23,
        64'hfc043783_fcf43823,
        64'hfc843783_fef43023,
        64'hfd878793_03040793,
        64'h03143423_03043023,
        64'hec1ce818_e414fac4,
        64'h3c23fcb4_3023fca4,
        64'h34230880_e0a2e486,
        64'h71198082_61457402,
        64'h70a2853e_87aab9ef,
        64'hf0efbf65_0513ffff,
        64'hf517fe84_3583fe04,
        64'h3603fd84_3683fd04,
        64'h3703fcd4_3823fcc4,
        64'h3c23feb4_3023fea4,
        64'h34231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_87aabdef,
        64'hf0efc945_0513ffff,
        64'hf51785be_567dfd84,
        64'h3683fd04_3703fe84,
        64'h0793fcb4_3823fca4,
        64'h3c231800_f022f406,
        64'h71798082_61657442,
        64'h70e2853e_fec42783,
        64'hfef42623_87aac1ef,
        64'hf0efc765_0513ffff,
        64'hf517fd84_3583fd04,
        64'h3603fc84_3683873e,
        64'hfe043783_fef43023,
        64'hfd878793_03040793,
        64'h03143423_03043023,
        64'hec1ce818_e414fcc4,
        64'h3423fcb4_3823fca4,
        64'h3c230080_f822fc06,
        64'h71598082_61257402,
        64'h70a2853e_fec42783,
        64'hfef42623_87aac7ef,
        64'hf0efcd65_0513ffff,
        64'hf517fd84_3583567d,
        64'hfd043683_873efe04,
        64'h3783fef4_3023fd07,
        64'h87930304_07930314,
        64'h34230304_3023ec1c,
        64'he818e414_e010fcb4,
        64'h3823fca4_3c231800,
        64'hf022f406_711d8082,
        64'h61097442_70e2853e,
        64'hfec42783_fef42623,
        64'h87aacdaf_f0efd905,
        64'h0513ffff_f51785be,
        64'h567dfc84_3683fd84,
        64'h0793fe04_3703fef4,
        64'h3023fc87_87930404,
        64'h07930314_3c230304,
        64'h3823f41c_f018ec14,
        64'he810e40c_fca43423,
        64'h0080f822_fc067119,
        64'h8082610d_644a60ea,
        64'h853e2781_fd843783,
        64'h97024501_f9043583,
        64'h863ef884_3683f984,
        64'h3703fd84_3783a019,
        64'h17fdf884_378300f7,
        64'h6663f884_3783fd84,
        64'h3703d807_99630007,
        64'hc783f804_37830001,
        64'hf8f43023_0785f804,
        64'h37839702_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_37830007,
        64'hc503f804_3783a80d,
        64'hf8f43023_0785f804,
        64'h37839702_02500513,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h3783a8b9_f8f43023,
        64'h0785f804_3783fca4,
        64'h3c23ba2f_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_36838736,
        64'h47814841_88bae03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_270386be,
        64'h639cf6e4_3c230087,
        64'h8713f784_3783a089,
        64'hfca43c23_cfcff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h87364781_484188ba,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442703,
        64'h86be639c_f6e43c23,
        64'h00878713_f7843783,
        64'hc3b10ff7_f793fbb4,
        64'h4783faf4_0da34785,
        64'hfef42623_0217e793,
        64'hfec42783_fef42423,
        64'h47c1a239_f8f43023,
        64'h0785f804_3783fce7,
        64'he7e32701_fe842703,
        64'hfce42223_0017871b,
        64'hfc442783_97020200,
        64'h0513f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_a00dcf8d,
        64'h27818b89_fec42783,
        64'hfbcdfee4_2223fff7,
        64'h871bfe44_2783d3e1,
        64'h27814007_f793fec4,
        64'h2783cf91_0007c783,
        64'hfc843783_9702f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'h0007c503_fce43423,
        64'h00178713_fc843783,
        64'ha03dfce7_e7e32701,
        64'hfe842703_fce42223,
        64'h0017871b_fc442783,
        64'h97020200_0513f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'ha00de7a5_27818b89,
        64'hfec42783_fcf42223,
        64'h87b200d7_73630006,
        64'h071b0007_869bfe44,
        64'h2783fc44_2603cf91,
        64'h27814007_f793fec4,
        64'h2783fcf4_222387aa,
        64'h8aaff0ef_fc843503,
        64'h85be57fd_a011fe44,
        64'h6783c781_2781fe44,
        64'h2783fcf4_3423639c,
        64'hf6e43c23_00878713,
        64'hf7843783_a4a1f8f4,
        64'h30230785_f8043783,
        64'hfce7e7e3_2701fe84,
        64'h2703fce4_28230017,
        64'h871bfd04_27839702,
        64'h02000513_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_3783a00d,
        64'hcf8d2781_8b89fec4,
        64'h27839702_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_37830ff7,
        64'hf513439c_f6e43c23,
        64'h00878713_f7843783,
        64'hfce7e7e3_2701fe84,
        64'h2703fce4_28230017,
        64'h871bfd04_27839702,
        64'h02000513_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_3783a00d,
        64'hef8d2781_8b89fec4,
        64'h2783fcf4_28234785,
        64'ha631f8f4_30230785,
        64'hf8043783_fca43c23,
        64'he50ff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_47818836,
        64'h88b2e03e_fe842783,
        64'he43efec4_2783fe44,
        64'h2603fd44_6683fb44,
        64'h6703faf4_2a232781,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783a801,
        64'h278193c1_17c2439c,
        64'hf6e43c23_00878713,
        64'hf7843783_cf812781,
        64'h0807f793_fec42783,
        64'ha8152781_0ff7f793,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783cf81,
        64'h27810407_f793fec4,
        64'h2783a841_fca43c23,
        64'hee0ff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_47818836,
        64'h88b2e03e_fe842783,
        64'he43efec4_2783fe44,
        64'h2603fd44_66836398,
        64'hf6e43c23_00878713,
        64'hf7843783_c3b12781,
        64'h1007f793_fec42783,
        64'ha8f9fca4_3c23847f,
        64'hf0eff984_3503f904,
        64'h3583fd84_3603f884,
        64'h36834781_883688b2,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442603,
        64'hfd446683_6398f6e4,
        64'h3c230087_8713f784,
        64'h3783c3b1_27812007,
        64'hf793fec4_2783a235,
        64'hfca43c23_f7cff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h87b68832_88aee03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_2583fd44,
        64'h66030ff7_f69301f7,
        64'hd79bfb04_27839301,
        64'h02079713_27812781,
        64'h40f707bb_8f3dfb04,
        64'h270341f7_d79bfb04,
        64'h2783faf4_2823439c,
        64'hf6e43c23_00878713,
        64'hf7843783_a8012781,
        64'h4107d79b_0107979b,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783cf91,
        64'h27810807_f793fec4,
        64'h2783a81d_27810ff7,
        64'hf793439c_f6e43c23,
        64'h00878713_f7843783,
        64'hcf812781_0407f793,
        64'hfec42783_a2cdfca4,
        64'h3c23833f_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_3683872e,
        64'h87ba8836_88b2e03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_2603fd44,
        64'h66830ff7_f71393fd,
        64'hfa843783_85be8f99,
        64'h8fb9fa84_378343f7,
        64'hd713fa84_3783faf4,
        64'h3423639c_f6e43c23,
        64'h00878713_f7843783,
        64'hc3bd2781_1007f793,
        64'hfec42783_ac89fca4,
        64'h3c239bbf_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_3683872e,
        64'h87ba8836_88b2e03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_2603fd44,
        64'h66830ff7_f71393fd,
        64'hfa043783_85be8f99,
        64'h8fb9fa04_378343f7,
        64'hd713fa04_3783faf4,
        64'h3023639c_f6e43c23,
        64'h00878713_f7843783,
        64'hc3bd2781_2007f793,
        64'hfec42783_18f71d63,
        64'h06400793_873e0007,
        64'hc783f804_378300f7,
        64'h0b630690_0793873e,
        64'h0007c783_f8043783,
        64'hfef42623_9bf9fec4,
        64'h2783c791_27814007,
        64'hf793fec4_2783fef4,
        64'h26239bcd_fec42783,
        64'h00f70763_06400793,
        64'h873e0007_c783f804,
        64'h378302f7_00630690,
        64'h0793873e_0007c783,
        64'hf8043783_fef42623,
        64'h0207e793_fec42783,
        64'h00f71863_05800793,
        64'h873e0007_c783f804,
        64'h3783fef4_26239bbd,
        64'hfec42783_fcf42a23,
        64'h47a9a809_fcf42a23,
        64'h478900f7_16630620,
        64'h0793873e_0007c783,
        64'hf8043783_a035fcf4,
        64'h2a2347a1_00f71663,
        64'h06f00793_873e0007,
        64'hc783f804_3783a099,
        64'hfcf42a23_47c100f7,
        64'h16630580_0793873e,
        64'h0007c783_f8043783,
        64'h00f70b63_07800793,
        64'h873e0007_c783f804,
        64'h37838782_97bad467,
        64'h87930000_57970007,
        64'h871b439c_97bad567,
        64'h87930000_57970027,
        64'h97139381_02069793,
        64'h6ce7e363_05300793,
        64'h0006871b_fdb7869b,
        64'h27810007_c783f804,
        64'h37830001_a0110001,
        64'ha0210001_a031f8f4,
        64'h30230785_f8043783,
        64'hfef42623_1007e793,
        64'hfec42783_a015f8f4,
        64'h30230785_f8043783,
        64'hfef42623_1007e793,
        64'hfec42783_a835f8f4,
        64'h30230785_f8043783,
        64'hfef42623_1007e793,
        64'hfec42783_a889f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0407e793,
        64'hfec42783_06f71663,
        64'h06800793_873e0007,
        64'hc783f804_3783f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0807e793,
        64'hfec42783_a079f8f4,
        64'h30230785_f8043783,
        64'hfef42623_2007e793,
        64'hfec42783_0af71463,
        64'h06c00793_873e0007,
        64'hc783f804_3783f8f4,
        64'h30230785_f8043783,
        64'hfef42623_1007e793,
        64'hfec42783_878297ba,
        64'he0c78793_00005797,
        64'h0007871b_439c97ba,
        64'he1c78793_00005797,
        64'h00279713_93810206,
        64'h97930ee7_e96347c9,
        64'h0006871b_f987869b,
        64'h27810007_c783f804,
        64'h3783f8f4_30230785,
        64'hf8043783_fef42223,
        64'h27814781_00075363,
        64'h0007871b_fbc42783,
        64'hfaf42e23_439cf6e4,
        64'h3c230087_8713f784,
        64'h378302f7_1a6302a0,
        64'h0793873e_0007c783,
        64'hf8043783_a091fef4,
        64'h222387aa_f86ff0ef,
        64'h853ef804_0793cb91,
        64'h87aaf54f_f0ef853e,
        64'h0007c783_f8043783,
        64'hf8f43023_0785f804,
        64'h3783fef4_26234007,
        64'he793fec4_278308f7,
        64'h106302e0_0793873e,
        64'h0007c783_f8043783,
        64'hfe042223_f8f43023,
        64'h0785f804_3783fef4,
        64'h2423fc04_2783a029,
        64'hfef42423_278140f0,
        64'h07bbfc04_2783fef4,
        64'h26230027_e793fec4,
        64'h27830207_d0632781,
        64'hfc042783_fcf42023,
        64'h439cf6e4_3c230087,
        64'h8713f784_378304f7,
        64'h176302a0_0793873e,
        64'h0007c783_f8043783,
        64'ha8b9fef4_242387aa,
        64'h833ff0ef_853ef804,
        64'h0793cb91_87aa801f,
        64'hf0ef853e_0007c783,
        64'hf8043783_fe042423,
        64'hf3852781_fe042783,
        64'h0001fe04_2023a021,
        64'hfef42023_4785f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0107e793,
        64'hfec42783_a01dfef4,
        64'h20234785_f8f43023,
        64'h0785f804_3783fef4,
        64'h26230087_e793fec4,
        64'h2783a091_fef42023,
        64'h4785f8f4_30230785,
        64'hf8043783_fef42623,
        64'h0047e793_fec42783,
        64'ha08dfef4_20234785,
        64'hf8f43023_0785f804,
        64'h3783fef4_26230027,
        64'he793fec4_2783a041,
        64'hfef42023_4785f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0017e793,
        64'hfec42783_878297ba,
        64'hfc078793_00005797,
        64'h0007871b_439c97ba,
        64'hfd078793_00005797,
        64'h00279713_93810206,
        64'h97930ce7_e06347c1,
        64'h0006871b_fe07869b,
        64'h27810007_c783f804,
        64'h3783fe04_2623f8f4,
        64'h30230785_f8043783,
        64'h2270006f_f8f43023,
        64'h0785f804_37839702,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h37830007_c503f804,
        64'h378302f7_0b630250,
        64'h0793873e_0007c783,
        64'hf8043783_26b0006f,
        64'hf8f43c23_86678793,
        64'h00000797_26079de3,
        64'hf9043783_fc043c23,
        64'hf6e43c23_f8d43023,
        64'hf8c43423_f8b43823,
        64'hf8a43c23_1100e922,
        64'hed067135_8082610d,
        64'h644a60ea_853e87aa,
        64'hb47ff0ef_fb843503,
        64'hfb043583_fa843603,
        64'hfa043683_fe843783,
        64'h883688b2_e03ef904,
        64'h2783e43e_401ce83e,
        64'h441cfc04_0713f974,
        64'h46830007_861bf884,
        64'h3783f6e7_ffe347fd,
        64'hfe843703_c791f984,
        64'h3783f8f4_3c2302f7,
        64'h57b3f884_3783f984,
        64'h3703fcf7_08239736,
        64'hff040693_fed43423,
        64'h00170693_fe843703,
        64'h0ff7f793_37d90ff7,
        64'hf7939fb9_fe744703,
        64'h06100793_a0190410,
        64'h0793c781_27810207,
        64'hf793441c_a01d0ff7,
        64'hf7930307_879bfe74,
        64'h478300e7_e96347a5,
        64'h0ff7f713_fe744783,
        64'hfef403a3_02f777b3,
        64'hf8843783_f9843703,
        64'hc7c1f984_3783c781,
        64'h27814007_f793441c,
        64'hc41c9bbd_441ce781,
        64'hf9843783_fe043423,
        64'hf8f42823_87baf8f4,
        64'h0ba38746_f9043423,
        64'hf8e43c23_fad43023,
        64'hfac43423_fab43823,
        64'hfaa43c23_1100e922,
        64'hed067135_8082610d,
        64'h644a60ea_853e87aa,
        64'hc5fff0ef_fb843503,
        64'hfb043583_fa843603,
        64'hfa043683_fe843783,
        64'h883688b2_e03ef904,
        64'h2783e43e_401ce83e,
        64'h441cfc04_0713f974,
        64'h46830007_861bf884,
        64'h3783f6e7_ffe347fd,
        64'hfe843703_c791f984,
        64'h3783f8f4_3c2302f7,
        64'h57b3f884_3783f984,
        64'h3703fcf7_08239736,
        64'hff040693_fed43423,
        64'h00170693_fe843703,
        64'h0ff7f793_37d90ff7,
        64'hf7939fb9_fe744703,
        64'h06100793_a0190410,
        64'h0793c781_27810207,
        64'hf793441c_a01d0ff7,
        64'hf7930307_879bfe74,
        64'h478300e7_e96347a5,
        64'h0ff7f713_fe744783,
        64'hfef403a3_02f777b3,
        64'hf8843783_f9843703,
        64'hc7c1f984_3783c781,
        64'h27814007_f793441c,
        64'hc41c9bbd_441ce781,
        64'hf9843783_fe043423,
        64'hf8f42823_87baf8f4,
        64'h0ba38746_f9043423,
        64'hf8e43c23_fad43023,
        64'hfac43423_fab43823,
        64'hfaa43c23_1100e922,
        64'hed067135_80826161,
        64'h640660a6_853e87aa,
        64'hc65ff0ef_fe843503,
        64'hfe043583_fd843603,
        64'hfd043683_fc843703,
        64'hfc043783_883e88ba,
        64'h441c4818_00e78023,
        64'h02000713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_3783cf91,
        64'h27818ba1_481ca015,
        64'h00e78023_02b00713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h3783cf99_27818b91,
        64'h481ca0a1_00e78023,
        64'h02d00713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_3783cf99,
        64'h0ff7f793_fbf44783,
        64'h06e7e863_47fdfc04,
        64'h370300e7_80230300,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_00e7ef63,
        64'h47fdfc04_370300e7,
        64'h80230620_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'h00e7ef63_47fdfc04,
        64'h370302f7_14634789,
        64'h0007871b_fb842783,
        64'ha81500e7_80230580,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_02e7e063,
        64'h47fdfc04_3703c785,
        64'h27810207_f793481c,
        64'h02f71a63_47c10007,
        64'h871bfb84_2783a88d,
        64'h00e78023_07800713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h378302e7_e06347fd,
        64'hfc043703_e7852781,
        64'h0207f793_481c02f7,
        64'h1a6347c1_0007871b,
        64'hfb842783_fcf43023,
        64'h17fdfc04_378300f7,
        64'h176347c1_0007871b,
        64'hfb842783_cf89fc04,
        64'h3783fcf4_302317fd,
        64'hfc043783_02f71663,
        64'hfc043703_00846783,
        64'h00f70863_fc043703,
        64'h00046783_c3a9fc04,
        64'h3783e7a1_27814007,
        64'hf793481c_12078363,
        64'h27818bc1_481cfce7,
        64'hf6e347fd_fc043703,
        64'h00f77763_fc043703,
        64'h00846783_cf812781,
        64'h8b85481c_00e78023,
        64'h03000713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_3783a831,
        64'hfce7fae3_47fdfc04,
        64'h370302f7_7563fc04,
        64'h37030004_678300e7,
        64'h80230300_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'ha831c41c_37fd441c,
        64'hc3952781_8bb1481c,
        64'he7890ff7_f793fbf4,
        64'h4783cb9d_27818b85,
        64'h481ccf9d_2781441c,
        64'hebd12781_8b89481c,
        64'hfaf42c23_87bafaf4,
        64'h0fa38746_87c2fcf4,
        64'h3023fce4_3423fcd4,
        64'h3823fcc4_3c23feb4,
        64'h3023fea4_34230880,
        64'he0a2e486_715d8082,
        64'h61256446_60e6853e,
        64'hfc843783_fcf769e3,
        64'hfac46783_8f1dfe04,
        64'h3783fc84_37039702,
        64'h02000513_fd043583,
        64'h863efc04_3683fd84,
        64'h3703fce4_34230017,
        64'h8713fc84_3783a00d,
        64'hcb9d2781_8b89fa84,
        64'h2783f7e1_fb043783,
        64'h9702fd04_3583863e,
        64'hfc043683_fd843703,
        64'hfce43423_00178713,
        64'hfc843783_0007c503,
        64'h97bafb04_3783fb84,
        64'h3703faf4_382317fd,
        64'hfb043783_a81dfcf7,
        64'h67e3fe84_3703fac4,
        64'h6783fef4_34230785,
        64'hfe843783_97020200,
        64'h0513fd04_3583863e,
        64'hfc043683_fd843703,
        64'hfce43423_00178713,
        64'hfc843783_a035fef4,
        64'h3423fb04_3783efa5,
        64'h27818b85_fa842783,
        64'he3c92781_8b89fa84,
        64'h2783fef4_3023fc84,
        64'h3783faf4_242387ba,
        64'hfaf42623_874687c2,
        64'hfaf43823_fae43c23,
        64'hfcd43023_fcc43423,
        64'hfcb43823_fca43c23,
        64'h1080e8a2_ec86711d,
        64'h80826145_740270a2,
        64'h853efec4_2783ffc5,
        64'h87aaf6df_f0ef853e,
        64'h0007c783_639cfd84,
        64'h3783fef4_2623fd07,
        64'h879b2781_9fb92781,
        64'h0007c783_e290fd84,
        64'h36830017_8613639c,
        64'hfd843783_0007871b,
        64'h0017979b_9fb90027,
        64'h979b87ba_fec42703,
        64'ha825fe04_2623fca4,
        64'h3c231800_f022f406,
        64'h71798082_61056462,
        64'h853e0ff7_f7938b85,
        64'h4781a011_478500e7,
        64'he4630390_07930ff7,
        64'hf713fef4_478300e7,
        64'hfc6302f0_07930ff7,
        64'hf713fef4_4783fef4,
        64'h07a387aa_1000ec22,
        64'h11018082_61457422,
        64'h853e2781_40f707b3,
        64'hfd843783_fe843703,
        64'hf3e5fce4_3823fff7,
        64'h8713fd04_3783cb81,
        64'h0007c783_fe843783,
        64'hfef43423_0785fe84,
        64'h3783a031_fef43423,
        64'hfd843783_fcb43823,
        64'hfca43c23_1800f422,
        64'h71798082_61457402,
        64'h70a20001_9682853e,
        64'h85bafef4_47836798,
        64'hfe043783_6394fe04,
        64'h3783cf81_0ff7f793,
        64'hfef44783_fef407a3,
        64'hfcd43823_fcc43c23,
        64'hfeb43023_87aa1800,
        64'hf022f406_71798082,
        64'h61457402_70a20001,
        64'h8b7ff0ef_853efef4,
        64'h4783c791_0ff7f793,
        64'hfef44783_fef407a3,
        64'hfcd43823_fcc43c23,
        64'hfeb43023_87aa1800,
        64'hf022f406_71798082,
        64'h61457422_0001fef4,
        64'h07a3fcd4_3823fcc4,
        64'h3c23feb4_302387aa,
        64'h1800f422_71798082,
        64'h61457422_000100e7,
        64'h8023fef4_470397ba,
        64'hfd843783_fe043703,
        64'h00f77b63_fd043783,
        64'hfd843703_fef407a3,
        64'hfcd43823_fcc43c23,
        64'hfeb43023_87aa1800,
        64'hf4227179_8082610d,
        64'h690a64aa_644a60ea,
        64'hf6040113_853e8126,
        64'h814a4781_2b0010ef,
        64'h84850513_00006517,
        64'ha80157f9_2c0010ef,
        64'h5f050513_00005517,
        64'h85befac4_27832d20,
        64'h10ef5ea5_05130000,
        64'h5517c395_2781fac4,
        64'h2783faf4_262387aa,
        64'hb33ff0ef_f6843503,
        64'h85be863a_f6442703,
        64'h2781739c_f7843783,
        64'h304010ef_88450513,
        64'h00006517_f6f43c23,
        64'hf8043783_eae7d2e3,
        64'h478d0007_871bfd04,
        64'h2783fcf4_28232785,
        64'hfd042783_330010ef,
        64'h8a850513_00006517,
        64'hfce7d6e3_04700793,
        64'h0007871b_fdc42783,
        64'hfcf42e23_2785fdc4,
        64'h27833560_10ef8465,
        64'h05130000_651785be,
        64'h27810387_c78397ba,
        64'hfdc42783_f7043703,
        64'ha02dfc04_2e2337a0,
        64'h10ef8da5_05130000,
        64'h65173860_10ef8ce5,
        64'h05130000_651785be,
        64'h7b9cf704_378339a0,
        64'h10ef8ca5_05130000,
        64'h651785be_779cf704,
        64'h37833ae0_10ef8c65,
        64'h05130000_651785be,
        64'h739cf704_3783fce7,
        64'hd7e347bd_0007871b,
        64'hfd842783_fcf42c23,
        64'h2785fd84_27833da0,
        64'h10ef8ca5_05130000,
        64'h651785be_27810107,
        64'hc78397ba_fd842783,
        64'hf7043703_a02dfc04,
        64'h2c233fe0_10ef8f65,
        64'h05130000_6517fce7,
        64'hd7e347bd_0007871b,
        64'hfd442783_fcf42a23,
        64'h2785fd44_27834220,
        64'h10ef9125_05130000,
        64'h651785be_27810007,
        64'hc78397ba_fd442783,
        64'hf7043703_a02dfc04,
        64'h2a234460_10ef9165,
        64'h05130000_65174520,
        64'h10ef90a5_05130000,
        64'h651785be_fd042783,
        64'hf6f43823_97ba2701,
        64'h0077171b_fd042703,
        64'hf8043783_aa91fc04,
        64'h2823aac9_57f94820,
        64'h10ef91a5_05130000,
        64'h651785be_fac42783,
        64'h494010ef_7ac50513,
        64'h00005517_c3952781,
        64'hfac42783_faf42623,
        64'h87aacf5f_f0ef853a,
        64'h85be4605_278167bc,
        64'hf9043783_f8043703,
        64'hf8f43023_00078793,
        64'h878a40f1_01330792,
        64'h839107bd_f8e43423,
        64'h177d873e_fc043783,
        64'h4e4010ef_95c50513,
        64'h00006517_85be4bfc,
        64'hf9043783_4f8010ef,
        64'h95050513_00006517,
        64'h85be4bbc_f9043783,
        64'h50c010ef_93c50513,
        64'h00006517_85be67bc,
        64'hf9043783_520010ef,
        64'h93850513_00006517,
        64'h85be739c_f9043783,
        64'h534010ef_93450513,
        64'h00006517_85be6f9c,
        64'hf9043783_548010ef,
        64'h93050513_00006517,
        64'h85be4bdc_f9043783,
        64'h55c010ef_92c50513,
        64'h00006517_85be4b9c,
        64'hf9043783_570010ef,
        64'h92850513_00006517,
        64'h85be47dc_f9043783,
        64'h584010ef_92450513,
        64'h00006517_85be479c,
        64'hf9043783_598010ef,
        64'h92050513_00006517,
        64'h85be639c_f9043783,
        64'h5ac010ef_91450513,
        64'h00006517_f8f43823,
        64'hf9843783_ae1157f9,
        64'h5c4010ef_8f450513,
        64'h00006517_85befac4,
        64'h27835d60_10ef8ee5,
        64'h05130000_6517c395,
        64'h2781fac4_2783faf4,
        64'h262387aa_e37ff0ef,
        64'h853e4585_4605f984,
        64'h3783f8f4_3c230007,
        64'h8793878a_40f10133,
        64'h07928391_07bdfae4,
        64'h3023177d_873e893a,
        64'h870afc04_3783f6e7,
        64'hefe3fc04_3703fcc4,
        64'h2783fcf4_26232791,
        64'hfcc42783_638010ef,
        64'h98850513_00006517,
        64'h873e2781_0ff7f793,
        64'h0007c783_97bafb04,
        64'h37032781_278dfcc4,
        64'h27830007_869b0ff7,
        64'hf7930007_c78397ba,
        64'hfb043703_27812789,
        64'hfcc42783_0007861b,
        64'h0ff7f793_0007c783,
        64'h97bafb04_37032781,
        64'h2785fcc4_27830007,
        64'h859b0ff7_f7930007,
        64'hc78397ba_fcc42783,
        64'hfb043703_a8b5fc04,
        64'h2623a111_57f96b20,
        64'h10ef9e25_05130000,
        64'h651785be_fac42783,
        64'h6c4010ef_9dc50513,
        64'h00006517_c3952781,
        64'hfac42783_faf42623,
        64'h87aaf25f_f0ef853e,
        64'h45854605_fb043783,
        64'hfaf43823_00078793,
        64'h878a40f1_01330792,
        64'h839107bd_fae43c23,
        64'h177d873e_fc043783,
        64'hfcf43023_20000793,
        64'h714010ef_a1450513,
        64'h00006517_a99d57fd,
        64'h724010ef_9fc50513,
        64'h00006517_cb892781,
        64'hfc842783_fcf42423,
        64'h87aaecdf_f0ef84be,
        64'h878af6f4_222387ae,
        64'hf6a43423_1100e14a,
        64'he526e922_ed067135,
        64'h80826145_740270a2,
        64'h853e4781_a01157fd,
        64'h76c010ef_a2450513,
        64'h00006517_85befec4,
        64'h2783cf81_2781fec4,
        64'h2783fef4_262387aa,
        64'h05b030ef_c3c50513,
        64'h1fff0517_85be4605,
        64'hfd843683_fd442783,
        64'hfcf42823_87bafcf4,
        64'h2a238732_87aefca4,
        64'h3c231800_f022f406,
        64'h71798082_61056442,
        64'h60e2853e_47817ca0,
        64'h10efa625_05130000,
        64'h6517a801_57f57da0,
        64'h10efa425_05130000,
        64'h651785be_fe442783,
        64'hcf812781_fe442783,
        64'hfef42223_87aa5900,
        64'h20efcaa5_05131fff,
        64'h0517a081_57f900b0,
        64'h10efa4a5_05130000,
        64'h651785be_fe442783,
        64'hcf812781_fe442783,
        64'hfef42223_87aa4db0,
        64'h10efcda5_05131fff,
        64'h0517fe84_3583863e,
        64'h43dcfe84_3783a8b5,
        64'h57fd0470_10efa665,
        64'h05130000_6517eb89,
        64'hfe843783_fea43423,
        64'h2b9010ef_45010630,
        64'h10efa6a5_05130000,
        64'h65171000_e822ec06,
        64'h11018082_61457402,
        64'h70a20001_eb9ff0ef,
        64'h01078513_07fa478d,
        64'h02000593_ec9ff0ef,
        64'h00878513_07fa478d,
        64'h0c700593_ed9ff0ef,
        64'h00c78513_07fa478d,
        64'h458dee7f_f0ef0047,
        64'h851307fa_478d85be,
        64'h0ff7f793_27810087,
        64'hd79bfec4_2783f03f,
        64'hf0ef01e7_9513478d,
        64'h85be0ff7_f793fec4,
        64'h2783f17f_f0ef00c7,
        64'h851307fa_478d0800,
        64'h0593f27f_f0ef0047,
        64'h851307fa_478d4581,
        64'hfef42623_02f757bb,
        64'hfdc42703_27810047,
        64'h979bfd84_2783fcf4,
        64'h2c2387ba_fcf42e23,
        64'h872e87aa_1800f022,
        64'hf4067179_80826105,
        64'h644260e2_0001f6bf,
        64'hf0ef01e7_9513478d,
        64'h85befef4_4783dfed,
        64'h87aafc9f_f0ef0001,
        64'hfef407a3_87aa1000,
        64'he822ec06_11018082,
        64'h01416402_60a2853e,
        64'h27810207_f7932781,
        64'h87aafd3f_f0ef0147,
        64'h851307fa_478d0800,
        64'he022e406_11418082,
        64'h61056462_853e0ff7,
        64'hf7930007_c783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826145,
        64'h74220001_00e78023,
        64'hfd744703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf40ba3_87aefca4,
        64'h3c231800_f4227179,
        64'ha0011cf0_10efbae5,
        64'h05130000_65178402,
        64'h19858593_00006597,
        64'h10000437_eb812781,
        64'hfe842783_fef42423,
        64'h87aa29e0_00ef1000,
        64'h053765a1_fce7dae3,
        64'h47910007_871bfec4,
        64'h2783fef4_26232785,
        64'hfec42783_219010ef,
        64'hbf050513_00006517,
        64'h437010ef_24078513,
        64'h000f47b7_a015fe04,
        64'h26232370_10efbe65,
        64'h05130000_651711e0,
        64'h00efa007_85130262,
        64'h67b72007_859367f1,
        64'h1000e822_ec061101,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00048067,
        64'h100004b7_29458593,
        64'h00006597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h0e4000ef_fec10113,
        64'h3fff0117_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
