/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 3529;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd0080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h08090000_38000000,
        64'hda0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'hffffb340_ffffb9dc,
        64'hffffb9dc_ffffb340,
        64'hffffb9dc_ffffb7c6,
        64'hffffb9dc_ffffb9dc,
        64'hffffb900_ffffb340,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb340,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb340_ffffb702,
        64'hffffb340_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb340_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9dc,
        64'hffffb9dc_ffffb9b0,
        64'hffffb32a_ffffb342,
        64'hffffb342_ffffb342,
        64'hffffb342_ffffb342,
        64'hffffb2fa_ffffb342,
        64'hffffb342_ffffb342,
        64'hffffb342_ffffb342,
        64'hffffb342_ffffb342,
        64'hffffb27a_ffffb342,
        64'hffffb312_ffffb342,
        64'hffffb2ba_ffffb0c6,
        64'hffffb15c_ffffb15c,
        64'hffffb0e4_ffffb15c,
        64'hffffb102_ffffb15c,
        64'hffffb15c_ffffb15c,
        64'hffffb15c_ffffb15c,
        64'hffffb15c_ffffb15c,
        64'hffffb13e_ffffb15c,
        64'hffffb15c_ffffb120,
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00586c6c_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000000_00007525,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000000_00007525,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_58323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h000a5838_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h000a5838_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_000a586c,
        64'h6c363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h00000000_0a756c6c,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h00000000_0a756c6c,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_0a583830,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_0a583830,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_0a583830,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_0a583830,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h00000000_0000000a,
        64'h00000000_00006325,
        64'h00202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h00000000_0a642520,
        64'h3a737574_61747320,
        64'h2c64656c_69616620,
        64'h64616552_20304453,
        64'h00000000_0a216465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a6425,
        64'h203a7375_74617473,
        64'h202c6465_6c696166,
        64'h206e6f69_74617a69,
        64'h6c616974_696e6920,
        64'h64726163_20304453,
        64'h0000000a_6425203a,
        64'h73757461_7473202c,
        64'h64656c69_6166206c,
        64'h61697469_6e692067,
        64'h69666e6f_63204453,
        64'h00000000_0000000a,
        64'h2164656c_69616620,
        64'h6769666e_6f632070,
        64'h756b6f6f_6c204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_0000000a,
        64'h00000000_002e2e2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00008082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'h930fc0ef_4505a031,
        64'hfef42623_4785e789,
        64'h27810807_f7932781,
        64'h87aaa21f_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h37830001_a011f6e7,
        64'hfee30270_07930ff7,
        64'hf713fe94_4783fef4,
        64'h04a32785_fe944783,
        64'hcf992781_0407f793,
        64'h278187aa_a5bfe0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_a0adfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaa45f_d0effd84,
        64'h35035007_85936785,
        64'h46014685_a829fef4,
        64'h262387aa_a5ffd0ef,
        64'hfd843503_30078593,
        64'h67854601_468500f7,
        64'h1f634785_873e0347,
        64'hc783fd84_3783a8ad,
        64'hfe0404a3_9ecfc0ef,
        64'h4505b03f_e0ef853e,
        64'h03e00593_863afe64,
        64'h570343dc_fd843783,
        64'hfef41323_0407e793,
        64'hfe645783_fef41323,
        64'h87aaaf1f_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h37838ee7_92234741,
        64'h1ffeb797_b45fe0ef,
        64'h853e4591_863afea4,
        64'h570343dc_fd843783,
        64'hfef41523_8ff917fd,
        64'h6785fea4_5703fef4,
        64'h15230017_979bfea4,
        64'h5783aa35_478590e7,
        64'hae234705_1ffeb797,
        64'h85efc0ef_78c50513,
        64'h00000517_78458593,
        64'h00000597_4a200613,
        64'ha02502f7_1c63478d,
        64'h873e0377_c783fd84,
        64'h3783fef4_15230400,
        64'h07939407_ab231ffe,
        64'hb797a251_478596e7,
        64'ha2234705_1ffeb797,
        64'h8a6fc0ef_7d450513,
        64'h00000517_7cc58593,
        64'h00000597_4a100613,
        64'ha02504f7_17631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_37839807,
        64'had231ffe_b797c385,
        64'hfd843783_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aab7ff_e0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783c3ff,
        64'he0ef853e_03000593,
        64'h460943dc_fd843783,
        64'hdfc52781_8b89fe84,
        64'h2783a83d_fef42623,
        64'h4785c63f_e0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hc3852781_8ff967a1,
        64'hfe842703_fef42423,
        64'h87aac51f_e0ef853e,
        64'h03000593_43dcfd84,
        64'h3783a8bd_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hc3bfd0ef_fd843503,
        64'h60000593_863e4681,
        64'hfd442783_fcf42a23,
        64'h87aefca4_3c231800,
        64'hf022f406_71798082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'hc45fe0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfc843783_d05fe0ef,
        64'h853e0300_05934609,
        64'h43dcfc84_3783dfc5,
        64'h27818b89_fdc42783,
        64'ha83dfef4_26234785,
        64'hd29fe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fc84_3783c385,
        64'h27818ff9_67a1fdc4,
        64'h2703fcf4_2e2387aa,
        64'hd17fe0ef_853e0300,
        64'h059343dc_fc843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aad01f,
        64'hd0effc84_35038007,
        64'h85936785_863e4685,
        64'hfe442783_b2e79b23,
        64'h47451ffe_b7970ff0,
        64'h000ff46f_e0effc84,
        64'h350385be_fc043603,
        64'h2781fe24_5783daff,
        64'he0ef853e_4591863a,
        64'hfe045703_43dcfc84,
        64'h3783fef4_10238ff9,
        64'h17fd6785_fe045703,
        64'hfef41023_20000793,
        64'hfef41123_4785fce7,
        64'hdee31ff0_07930007,
        64'h871bfe84_2783fef4,
        64'h24232785_fe842783,
        64'h00078023_97bafc04,
        64'h3703fe84_2783a225,
        64'h4785bae7_a8234705,
        64'h1ffeb797_af2fc0ef,
        64'ha2050513_00001517,
        64'ha1858593_00001597,
        64'h36900613_a081fe04,
        64'h2423bc07_ab231ffe,
        64'hb797aab1_4785bee7,
        64'ha2234705_1ffeb797,
        64'hb26fc0ef_a5450513,
        64'h00001517_a4c58593,
        64'h00001597_36800613,
        64'ha02502f7_1d631117,
        64'h87931111_17b7873e,
        64'h53dcfc84_3783c007,
        64'had231ffe_b797c385,
        64'hfc843783_fe042223,
        64'hfcb43023_fca43423,
        64'h0080f822_fc067139,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623a019_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'he4bfd0ef_fd843503,
        64'ha0078593_67ad4601,
        64'h4681a03d_fef42623,
        64'h4785a82d_4785c8e7,
        64'ha2234705_1ffeb797,
        64'hbc6fc0ef_af450513,
        64'h00001517_aec58593,
        64'h00001597_33900613,
        64'ha025cb8d_2781fec4,
        64'h2783fef4_262387aa,
        64'he9bfd0ef_fd843503,
        64'h70078593_678d863e,
        64'h46814bbc_fd843783,
        64'hcc07a623_1ffeb797,
        64'ha8414785_cce7ad23,
        64'h47051ffe_b797c1cf,
        64'hc0efb4a5_05130000,
        64'h1517b425_85930000,
        64'h15973380_0613a025,
        64'h04f71e63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_d007a823,
        64'h1ffeb797_c385fd84,
        64'h3783fca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'hfe842783_fe042423,
        64'hf99fe0ef_853a02c0,
        64'h0593863e_93c117c2,
        64'h0047e793_fe445783,
        64'h43d8fd84_3783fef4,
        64'h122387aa_f83fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_d3e52781,
        64'h8b892781_fe645783,
        64'hfef41323_87aafa5f,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783a821,
        64'hfef41323_87aafbdf,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783806f,
        64'hf0ef853e_02c00593,
        64'h863afe44_570343dc,
        64'hfd843783_fef41223,
        64'h0017e793_93c117c2,
        64'h8fd9fe44_5783fec4,
        64'h5703fef4_1623f007,
        64'hf793fec4_5783fef4,
        64'h16230087_979bfec4,
        64'h5783fef4_12230ff7,
        64'hf793fe44_5783fef4,
        64'h122387aa_822ff0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a0a586ef,
        64'hf0ef853e_02c00593,
        64'h863afe44_570343dc,
        64'hfd843783_fef41223,
        64'h0017e793_93c117c2,
        64'h8fd9fe44_57839341,
        64'h03079713_8fd9fe24,
        64'h5783fec4_5703fef4,
        64'h1623f007_f793fec4,
        64'h5783fef4_16230087,
        64'h979bfec4_5783fef4,
        64'h11230c07_f793fe24,
        64'h5783fef4_11230067,
        64'h979bfe24_5783fef4,
        64'h11230087_d79bfec4,
        64'h5783fef4_122303f7,
        64'hf793fe44_5783fef4,
        64'h122387aa_8baff0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_08f71e63,
        64'h4789873e_0367c783,
        64'hfd843783_a249fef4,
        64'h24234785_00e7f663,
        64'h10000793_0007871b,
        64'hfee45783_fae7fee3,
        64'h10000793_0007871b,
        64'hfee45783_fef41723,
        64'h0017979b_fee45783,
        64'ha839fef4_16230017,
        64'hd79bfee4_578300e7,
        64'he9632781_fd442783,
        64'h0007871b_02f757bb,
        64'h2781fee4_57834798,
        64'hfd843783_a82dfef4,
        64'h17234785_a2edfef4,
        64'h24234785_06e7fa63,
        64'h7fe00793_0007871b,
        64'hfee45783_fae7ffe3,
        64'h7fe00793_0007871b,
        64'hfee45783_fef41723,
        64'h2785fee4_5783a831,
        64'hfef41623_0017d79b,
        64'hfee45783_00e7e963,
        64'h2781fd44_27830007,
        64'h871b02f7_57bb2781,
        64'hfee45783_4798fd84,
        64'h3783a825_fef41723,
        64'h4785ac91_4785f8e7,
        64'ha6234705_1ffeb797,
        64'hecefc0ef_dfc50513,
        64'h00001517_df458593,
        64'h00001597_2c400613,
        64'ha02508f7_19634789,
        64'h873e0367_c783fd84,
        64'h3783a1af_f0ef853e,
        64'h02c00593_863afe44,
        64'h570343dc_fd843783,
        64'hfef41223_9be9fe44,
        64'h5783fef4_122387aa,
        64'ha06ff0ef_853e02c0,
        64'h059343dc_fd843783,
        64'hfe07aa23_1ffeb797,
        64'ha4e94785_00e7a123,
        64'h47051ffe_b797f44f,
        64'hc0efe725_05130000,
        64'h1517e6a5_85930000,
        64'h15972c30_0613a025,
        64'h06f71e63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_0207ac23,
        64'h1ffeb797_c385fd84,
        64'h3783fe04_1623fcf4,
        64'h2a2387ae_fca43c23,
        64'h1800f022_f4067179,
        64'h80826165_740670a6,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aaa26f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcf984_3783b66f,
        64'hf0ef853e_02800593,
        64'h863a0ff7_7713fe44,
        64'h270343dc_f9843783,
        64'hfef42223_0047e793,
        64'hfe442783_fef42223,
        64'h87aab58f_f0ef853e,
        64'h02800593_43dcf984,
        64'h3783a13f_c0ef3e80,
        64'h0513a09d_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h734000ef_f9843503,
        64'h02f71163_479d873e,
        64'h57fcf984_3783a849,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_0b8000ef,
        64'hf9843503_85be5f9c,
        64'hf9843783_b7cff0ef,
        64'h853e0300_05934609,
        64'h43dcf984_3783dfc5,
        64'h27818b89_fe442783,
        64'ha8d1fef4_26234785,
        64'hba0ff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8f984_3783c385,
        64'h27818ff9_67a1fe44,
        64'h2703fef4_222387aa,
        64'hb8eff0ef_853e0300,
        64'h059343dc_f9843783,
        64'haa11fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aab78f,
        64'he0eff984_35036000,
        64'h0593863e_4681fe84,
        64'h2783df98_5007071b,
        64'h03197737_f9843783,
        64'hfef42423_1007879b,
        64'h03b907b7_a831df98,
        64'h5007071b_03197737,
        64'hf9843783_fef42423,
        64'h1007879b_03b907b7,
        64'h02f71063_4791873e,
        64'h57fcf984_3783a099,
        64'hdf982007_071b0beb,
        64'hc737f984_3783fef4,
        64'h24232007_879b03b9,
        64'h07b702f7_1063479d,
        64'h873e57fc_f9843783,
        64'ha275fef4_26234785,
        64'h14078963_2781fec4,
        64'h2783fef4_262387aa,
        64'h1d4000ef_f9843503,
        64'h50078593_031977b7,
        64'hdf985007_071b0319,
        64'h7737f984_3783ca6f,
        64'hf0ef853e_03000593,
        64'h460943dc_f9843783,
        64'hdfc52781_8b89fe44,
        64'h2783aafd_fef42623,
        64'h4785ccaf_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_f9843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aacb8f_f0ef853e,
        64'h03000593_43dcf984,
        64'h3783ac3d_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hca2fe0ef_f9843503,
        64'h60000593_863e4681,
        64'hfe842783_fef42423,
        64'h1007879b_03b907b7,
        64'h0cf71663_4789873e,
        64'h0347c783_f9843783,
        64'ha451fef4_26234785,
        64'h22078563_2781fec4,
        64'h2783fef4_262387aa,
        64'h2ac000ef_f9843503,
        64'h85be5f9c_f9843783,
        64'hdf980807_071b02fa,
        64'hf737f984_3783d7ef,
        64'hf0ef853e_03000593,
        64'h460943dc_f9843783,
        64'hdfc52781_8b89fe44,
        64'h2783acd9_fef42623,
        64'h4785da2f_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_f9843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aad90f_f0ef853e,
        64'h03000593_43dcf984,
        64'h3783ae19_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hd7afe0ef_f9843503,
        64'h60000593_863e4685,
        64'hfe842783_fef42423,
        64'h37c58100_07b73ae7,
        64'h9c234745_1ffeb797,
        64'h0ff0000f_fc9fe0ef,
        64'hf9843503_85be863a,
        64'hfa040713_2781fe24,
        64'h5783e32f_f0ef853e,
        64'h4591863a_fe045703,
        64'h43dcf984_3783fef4,
        64'h10238ff9_17fd6785,
        64'hfe045703_fef41023,
        64'h04000793_fef41123,
        64'h4785a64d_478540e7,
        64'ha6234705_1ffeb797,
        64'hb4ffc0ef_27c50513,
        64'h00001517_27458593,
        64'h00001597_1fc00613,
        64'ha02514f7_13634785,
        64'h873e0347_c783f984,
        64'h37834207_af231ffe,
        64'hb797a6cd_478544e7,
        64'ha6234705_1ffeb797,
        64'hb8ffc0ef_2bc50513,
        64'h00001517_2b458593,
        64'h00001597_1fb00613,
        64'ha02504f7_13631117,
        64'h87931111_17b7873e,
        64'h53dcf984_37834807,
        64'ha1231ffe_b797c385,
        64'hf9843783_fc043c23,
        64'hfc043823_fc043423,
        64'hfc043023_fa043c23,
        64'hfa043823_fa043423,
        64'hfa043023_f8a43c23,
        64'h1880f0a2_f4867159,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aae86f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfc84_3783f46f,
        64'hf0ef853e_03000593,
        64'h460943dc_fc843783,
        64'hdfc52781_8b89fdc4,
        64'h2783a83d_fef42623,
        64'h4785f6af_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fc843783,
        64'hc3852781_8ff967a1,
        64'hfdc42703_fcf42e23,
        64'h87aaf58f_f0ef853e,
        64'h03000593_43dcfc84,
        64'h3783a8bd_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hf42fe0ef_fc843503,
        64'h60000593_863e4685,
        64'hfe042783_0ff0000f,
        64'hfef42023_37c10100,
        64'h07b758e7_92234745,
        64'h1ffeb797_990ff0ef,
        64'hfc843503_85befc04,
        64'h36032781_fe645783,
        64'hff8ff0ef_853e4591,
        64'h863afe44_570343dc,
        64'hfc843783_fef41223,
        64'h8ff917fd_6785fe44,
        64'h5703fef4_12230400,
        64'h0793fef4_13234785,
        64'hfce7dee3_03f00793,
        64'h0007871b_fe842783,
        64'hfef42423_2785fe84,
        64'h27830007_802397ba,
        64'hfc043703_fe842783,
        64'haa054785_5ee7ad23,
        64'h47051ffe_b797d3df,
        64'hc0ef46a5_05130000,
        64'h15174625_85930000,
        64'h15971a40_0613a081,
        64'hfe042423_6207a023,
        64'h1ffeb797_a2954785,
        64'h62e7a723_47051ffe,
        64'hb797d71f_c0ef49e5,
        64'h05130000_15174965,
        64'h85930000_15971a30,
        64'h0613a025_02f71d63,
        64'h11178793_111117b7,
        64'h873e53dc_fc843783,
        64'h6607a223_1ffeb797,
        64'hc385fc84_3783fcb4,
        64'h3023fca4_34230080,
        64'hf822fc06_71398082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'h84dff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_90dff0ef,
        64'h853e03e0_0593863a,
        64'h93411742_fe842703,
        64'h43dcfd84_3783fef4,
        64'h24238fd9_fe842783,
        64'h57f8fd84_3783fef4,
        64'h24238ff9_17e167c1,
        64'hfe842703_fef42423,
        64'h87aa911f_f0ef853e,
        64'h03e00593_43dcfd84,
        64'h378304f7_19634791,
        64'h873e57fc_fd843783,
        64'h9e9ff0ef_853e0280,
        64'h0593863a_0ff77713,
        64'hfe842703_43dcfd84,
        64'h3783fef4_24230027,
        64'he793fe84_2783a039,
        64'hfef42423_0207e793,
        64'hfe842783_00f71963,
        64'h478d873e_0377c783,
        64'hfd843783_fef42423,
        64'h87aa9f9f_f0ef853e,
        64'h02800593_43dcfd84,
        64'h37838b2f_d0ef3e80,
        64'h05139cbf_f0ef853e,
        64'h03000593_460943dc,
        64'hfd843783_dfc52781,
        64'h8b89fe84_2783a8f5,
        64'hfef42623_47859eff,
        64'hf0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c3852781,
        64'h8ff967a1_fe842703,
        64'hfef42423_87aa9ddf,
        64'hf0ef853e_03000593,
        64'h43dcfd84_3783aa35,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_9c7fe0ef,
        64'hfd843503_60000593,
        64'h863e4681_fe442783,
        64'hfef42223_1007879b,
        64'h03b707b7_a039fef4,
        64'h22235007_879b03b7,
        64'h07b700f7_19634791,
        64'h873e57fc_fd843783,
        64'ha02dfef4_22232007,
        64'h879b03b7_07b7a825,
        64'hfef42223_6007879b,
        64'h03b707b7_00f71963,
        64'h4791873e_57fcfd84,
        64'h378302f7_1763478d,
        64'h873e0377_c783fd84,
        64'h378302e7_8ba34709,
        64'hfd843783_a03102e7,
        64'h8ba3470d_fd843783,
        64'h00f71863_47a1873e,
        64'h4bdcfd84_378300f7,
        64'h1f634795_873e0347,
        64'hc783fd84_378302f7,
        64'h17634789_873e0367,
        64'hc783fd84_3783a431,
        64'hfef42623_47851207,
        64'h8c632781_fec42783,
        64'hfef42623_87aaa99f,
        64'he0effd84_35036007,
        64'h859367a1_863e4681,
        64'hfe442783_fef42223,
        64'h0377c783_fd843783,
        64'h02e78ba3_4709fd84,
        64'h3783ac81_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hadbfe0ef_fd843503,
        64'h70078593_678d863e,
        64'h46814bbc_fd843783,
        64'h06f71b63_4785873e,
        64'h0347c783_fd843783,
        64'ha479fe04_262300e7,
        64'he563478d_873e4bdc,
        64'hfd843783_a45d4785,
        64'h92e7ab23_47051ffe,
        64'hc797878f_d0ef7a65,
        64'h05130000_151779e5,
        64'h85930000_15971170,
        64'h0613a025_04f71063,
        64'h4789873e_0367c783,
        64'hfd843783_9607a423,
        64'h1ffec797_a4dd4785,
        64'h96e7ab23_47051ffe,
        64'hc7978b8f_d0ef7e65,
        64'h05130000_15177de5,
        64'h85930000_15971160,
        64'h0613a025_04f71363,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'h9a07a623_1ffec797,
        64'hc385fd84_3783fca4,
        64'h3c231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_b91ff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fd843783,
        64'hc51ff0ef_853e0300,
        64'h05934609_43dcfd84,
        64'h3783dfc5_27818b89,
        64'hfe042783_a83dfef4,
        64'h26234785_c75ff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c385_27818ff9,
        64'h67a1fe04_2703fef4,
        64'h202387aa_c63ff0ef,
        64'h853e0300_059343dc,
        64'hfd843783_a8bdfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aac4df_e0effd84,
        64'h35033007_859367ad,
        64'h460186be_2781fe64,
        64'h57830ff0_000fa8e7,
        64'h94234745_1ffec797,
        64'he94ff0ef_fd843503,
        64'h85befd04_36032781,
        64'hfe645783_cfdff0ef,
        64'h853e4591_863afe44,
        64'h570343dc_fd843783,
        64'hfef41223_8ff917fd,
        64'h6785fe44_5703fef4,
        64'h122347a1_fef41323,
        64'h4785a8f5_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hccbfe0ef_fd843503,
        64'h70078593_678d863e,
        64'h46814bbc_fd843783,
        64'hfce7dfe3_479d0007,
        64'h871bfe84_2783fef4,
        64'h24232785_fe842783,
        64'h00078023_97bafd04,
        64'h3703fe84_2783aa91,
        64'h4785b2e7_a4234705,
        64'h1ffec797_a6afd0ef,
        64'h99850513_00002517,
        64'h99058593_00002597,
        64'h0ba00613_a081fe04,
        64'h2423b407_a7231ffe,
        64'hc797a261_4785b4e7,
        64'hae234705_1ffec797,
        64'ha9efd0ef_9cc50513,
        64'h00002517_9c458593,
        64'h00002597_0b900613,
        64'ha02502f7_1d631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783b807,
        64'ha9231ffe_c797c385,
        64'hfd843783_fcb43823,
        64'hfca43c23_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623e1ff,
        64'hf0ef8536_4591863e,
        64'h93c117c2_8ff917fd,
        64'h6785fd64_570343d4,
        64'hfd843783_fef42623,
        64'h278187aa_d99ff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fd843783,
        64'ha081fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aadf9f,
        64'he0effd84_35036585,
        64'h863e4681_2781fd64,
        64'h5783a0ad_fef42623,
        64'h4785a89d_4785c2e7,
        64'haa234705_1ffec797,
        64'hb76fd0ef_aa450513,
        64'h00002517_a9c58593,
        64'h00002597_07f00613,
        64'ha025cb8d_27813037,
        64'hf793fe84_2783fef4,
        64'h242387aa_e19ff0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783c607_af231ffe,
        64'hc797a0f9_4785c8e7,
        64'ha6234705_1ffec797,
        64'hbcefd0ef_afc50513,
        64'h00002517_af458593,
        64'h00002597_07e00613,
        64'ha02504f7_1f631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783cc07,
        64'ha1231ffe_c797c385,
        64'hfd843783_fcf41b23,
        64'h87aefca4_3c231800,
        64'hf022f406_71798082,
        64'h61056442_60e20001,
        64'heb7ff0ef_853e85ba,
        64'hfea44703_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h052387ba_fef405a3,
        64'h87b6fef4_26238732,
        64'h86ae87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_853e87aa,
        64'hea9ff0ef_853e9381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef405a3_87bafef4,
        64'h2623872e_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e20001,
        64'hf63ff0ef_853e85ba,
        64'hfe845703_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h142387ba_fef405a3,
        64'h87b6fef4_26238732,
        64'h86ae87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_853e87aa,
        64'hf47ff0ef_853e9381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef405a3_87bafef4,
        64'h2623872e_87aa1000,
        64'he822ec06_11018082,
        64'h61457422_000100e7,
        64'h9023fd64_5703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_1b2387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61457422,
        64'h000100e7_8023fd74,
        64'h4703fe84_3783fef4,
        64'h3423fd84_3783fcf4,
        64'h0ba387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61056462_853e2781,
        64'h439cfe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826105_6462853e,
        64'h93c117c2_0007d783,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61056462_853e0ff7,
        64'hf7930007_c783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826161,
        64'h640660a6_853efec4,
        64'h2783fe04_2623d3f8,
        64'hfb843783_0007871b,
        64'h0097d79b_fd842783,
        64'hfcf42c23_02f707bb,
        64'hfe042783_fd842703,
        64'hfcf42c23_02f707bb,
        64'hfdc42703_27812785,
        64'hfd842783_fcf42c23,
        64'h8fd9fd84_27830007,
        64'h871b8ff9_c0078793,
        64'h6785873e_278100a7,
        64'h979bfd04_2783fcf4,
        64'h2c230167_d79bfcc4,
        64'h2783fcf4_2e232781,
        64'h00f717bb_47052781,
        64'h27892781_8b9d2781,
        64'h0077d79b_fcc42783,
        64'hfef42023_278100f7,
        64'h17bb4705_27818bbd,
        64'h27810087_d79bfd04,
        64'h278302e7_8aa3fb84,
        64'h37830ff7_f7138bbd,
        64'h0ff7f793_27810127,
        64'hd79bfd44_2783fcf4,
        64'h2a232781_87aa9b1f,
        64'hd0ef853e_93811782,
        64'h278127f1_43dcfb84,
        64'h3783fcf4_28232781,
        64'h87aa9cdf_d0ef853e,
        64'h93811782_278127e1,
        64'h43dcfb84_3783fcf4,
        64'h26232781_87aa9e9f,
        64'hd0ef853e_93811782,
        64'h278127d1_43dcfb84,
        64'h3783fcf4_24232781,
        64'h87aaa05f_d0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783a23d,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_9c6ff0ef,
        64'hfb843503_90078593,
        64'h6785863e_46814bbc,
        64'hfb843783_aab1fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa9f4f_f0effb84,
        64'h35033000_0593863e,
        64'h46814bbc_fb843783,
        64'hcbb81234_0737fb84,
        64'h3783c7f8_fb843783,
        64'h0007871b_87aab25f,
        64'hd0ef853e_45f143dc,
        64'hfb843783_c7b8fb84,
        64'h37830007_871b87aa,
        64'hb3ffd0ef_853e45e1,
        64'h43dcfb84_3783c3f8,
        64'hfb843783_0007871b,
        64'h87aab59f_d0ef853e,
        64'h45d143dc_fb843783,
        64'hc3b8fb84_37830007,
        64'h871b87aa_b73fd0ef,
        64'h853e45c1_43dcfb84,
        64'h3783aaed_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'ha92ff0ef_fb843503,
        64'h20000593_46014681,
        64'hdb984705_fb843783,
        64'hc7892781_8ff94000,
        64'h07b7fe84_2703fa07,
        64'hdde3fe84_2783fef4,
        64'h242387aa_b2ffd0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'haca1fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaaf0f,
        64'hf0effb84_35031000,
        64'h059340ff_86374681,
        64'ha091fe04_2423a459,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_b1eff0ef,
        64'hfb843503_45814601,
        64'h4681a46d_fef42623,
        64'h4785e789_27818ff9,
        64'h67c1fe44_2703fef4,
        64'h222387aa_baffd0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfb84,
        64'h3783cb8d_47dcfb84,
        64'h378302f7_0e634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfb843783_a6014785,
        64'h18e7af23_47051ffe,
        64'hc7978e1f_d0effee5,
        64'h05130000_2517fee5,
        64'h85930000_259767d0,
        64'h0613a025_04f71363,
        64'h4789873e_0367c783,
        64'hfb843783_1c07a823,
        64'h1ffec797_a6814785,
        64'h1ce7af23_47051ffe,
        64'hc797921f_d0ef02e5,
        64'h05130000_251702e5,
        64'h85930000_259767c0,
        64'h0613a025_04f71363,
        64'h11178793_111117b7,
        64'h873e53dc_fb843783,
        64'h2007aa23_1ffec797,
        64'hc385fb84_3783faa4,
        64'h3c230880_e0a2e486,
        64'h715d8082_61217442,
        64'h70e20001_0ff0000f,
        64'hcfdfd0ef_853a85be,
        64'h27810807_8793fd84,
        64'h37839301_02079713,
        64'h27810587_879b43dc,
        64'hfd843783_00e79123,
        64'h97b6078e_07c19381,
        64'h02061793_fd843683,
        64'h93410307_971302f7,
        64'h07bb0006_861b36fd,
        64'hfec42683_93c117c2,
        64'hfe442783_93410307,
        64'h9713fd44_278300e7,
        64'h90230230_071397ba,
        64'h078e07c1_93811782,
        64'hfd843703_278137fd,
        64'hfec42783_c3d897b6,
        64'h078e07c1_93810206,
        64'h1793fd84_36830007,
        64'h871b9fb9_0006861b,
        64'h36fdfec4_26832781,
        64'h0107979b_fe842783,
        64'h0007871b_fc843783,
        64'hf8e7ebe3_2781fe84,
        64'h27830007_871b37fd,
        64'hfec42783_fef42423,
        64'h2785fe84_27830007,
        64'h912397ba_078e07c1,
        64'hfe846783_fd843703,
        64'h00e79023_02100713,
        64'h97ba078e_07c1fe84,
        64'h6783fd84_3703c3d8,
        64'h97b6078e_07c1fe84,
        64'h6783fd84_36830007,
        64'h871b9fb9_27810107,
        64'h979bfe84_27830007,
        64'h871bfc84_3783a8b1,
        64'hfe042423_fef42623,
        64'h2785fec4_2783c791,
        64'h27818ff9_17fd67c1,
        64'h873e2781_02f707bb,
        64'hfe442783_fd442703,
        64'hfef42623_0107d79b,
        64'h278102f7_07bbfe44,
        64'h2783fd44_2703a835,
        64'hfef42623_478500f7,
        64'h766367c1_873e2781,
        64'h02f707bb_fe442783,
        64'hfd442703_fef42223,
        64'h8ff917fd_6785fe44,
        64'h2703fef4_222387aa,
        64'heb7fd0ef_853e4591,
        64'h43dcfd84_3783fe04,
        64'h2223fe04_2423fe04,
        64'h2623fcf4_2a23fcc4,
        64'h342387ae_fca43c23,
        64'h0080f822_fc067139,
        64'h80826145_740270a2,
        64'h853efec4_27830001,
        64'ha011fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aae08f,
        64'hf0effd84_35037000,
        64'h0593863e_46814bbc,
        64'hfd843783_fe042623,
        64'hfca43c23_1800f022,
        64'hf4067179_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623f7ff,
        64'hd0ef853e_03000593,
        64'h460943dc_fd843783,
        64'hdfc52781_8b89fe44,
        64'h2783a00d_fef42623,
        64'h4785fa3f_d0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aaf91f_d0ef853e,
        64'h03000593_43dcfd84,
        64'h3783a08d_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'heb2ff0ef_fd843503,
        64'h90078593_6789863e,
        64'h86bafd44_2783fd04,
        64'h27034ee7_97230270,
        64'h07131ffe_c797a879,
        64'hfef42623_4785c3b9,
        64'h2781fec4_2783fef4,
        64'h262387aa_eeeff0ef,
        64'hfd843503_80078593,
        64'h6789863e_86bafd44,
        64'h2783fd04_270352e7,
        64'h9423470d_1ffec797,
        64'h02f71f63_47850007,
        64'h871bfd04_27830ff0,
        64'h000f1460_00effd84,
        64'h350385be_fc843603,
        64'hfd042783_a8f5fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa0890_00effd84,
        64'h35032000_059302f7,
        64'h03632000_0793873e,
        64'h278187aa_fcffd0ef,
        64'h853e9381_17822781,
        64'h279143dc_fd843783,
        64'ha281fef4_26234785,
        64'he7892781_8ff967c1,
        64'hfe842703_fef42423,
        64'h87aaffdf_d0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'hcb8d47dc_fd843783,
        64'h02f70e63_400007b7,
        64'h873e2781_8ff9c000,
        64'h07b7873e_579cfd84,
        64'h378300f7_1f634789,
        64'h873e0367_c783fd84,
        64'h3783fcf4_282387ba,
        64'hfcf42a23_fcd43423,
        64'h873287ae_fca43c23,
        64'h0080f822_fc067139,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aa87cf_e0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783966f,
        64'he0ef853e_03000593,
        64'h460943dc_fd843783,
        64'hdfc52781_8b89fe44,
        64'h2783a83d_fef42623,
        64'h478598af_e0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aa978f_e0ef853e,
        64'h03000593_43dcfd84,
        64'h3783a8bd_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h89bff0ef_fd843503,
        64'h20078593_6785863e,
        64'h86bafd44_2783fd04,
        64'h27036ce7_9b230370,
        64'h07131ffe_c797a86d,
        64'hfef42623_4785c3b9,
        64'h2781fec4_2783fef4,
        64'h262387aa_8d7ff0ef,
        64'hfd843503_10078593,
        64'h6785863e_86bafd44,
        64'h2783fd04_270370e7,
        64'h9823474d_1ffec797,
        64'h02f71f63_47850007,
        64'h871bfd04_27830ff0,
        64'h000f32e0_00effd84,
        64'h350385be_fc843603,
        64'hfd042783_aa21fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa2710_00effd84,
        64'h35032000_059302f7,
        64'h03632000_0793873e,
        64'h278187aa_9b6fe0ef,
        64'h853e9381_17822781,
        64'h279143dc_fd843783,
        64'haab1fef4_26234785,
        64'he7892781_8ff967c1,
        64'hfe842703_fef42423,
        64'h87aa9e4f_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'hcb8d47dc_fd843783,
        64'h02f70e63_400007b7,
        64'h873e2781_8ff9c000,
        64'h07b7873e_579cfd84,
        64'h378300f7_1f634789,
        64'h873e0367_c783fd84,
        64'h3783fcf4_282387ba,
        64'hfcf42a23_fcd43423,
        64'h873287ae_fca43c23,
        64'h0080f822_fc067139,
        64'h80826145_7422853e,
        64'hfec42783_0001a011,
        64'h0001a021_0001a031,
        64'hfef42623_8fd9fd44,
        64'h2783fec4_2703a831,
        64'hfef42623_01a7e793,
        64'hfec42783_a02dfef4,
        64'h262303a7_e793fec4,
        64'h2783a825_fef42623,
        64'h01a7e793_fec42783,
        64'ha099fef4_26230027,
        64'he793fec4_2783a891,
        64'hfef42623_03a7e793,
        64'hfec42783_a08dfef4,
        64'h262303a7_e793fec4,
        64'h2783a885_fef42623,
        64'h01a7e793_fec42783,
        64'ha8bdfef4_26230097,
        64'he793fec4_2783a071,
        64'hfef42623_03a7e793,
        64'hfec42783_a869fef4,
        64'h262301a7_e793fec4,
        64'h278300f7_19634785,
        64'h873e0347_c783fd84,
        64'h3783a865_fef42623,
        64'h01a7e793_fec42783,
        64'ha0d9fef4_262301a7,
        64'he793fec4_2783a8d1,
        64'hfef42623_01b7e793,
        64'hfec42783_a0cdfef4,
        64'h262303a7_e793fec4,
        64'h278300f7_19634785,
        64'h873e0347_c783fd84,
        64'h3783a201_fef42623,
        64'h01b7e793_fec42783,
        64'ha239fef4_262301b7,
        64'he793fec4_2783aa31,
        64'hfef42623_0097e793,
        64'hfec42783_a22dfef4,
        64'h26230027_e793fec4,
        64'h2783aa39_0ef70563,
        64'h90078793_67ad0007,
        64'h871b10e6_8a633007,
        64'h0713672d_0007869b,
        64'h10e68a63_a0070713,
        64'h672d0007_869ba2a9,
        64'h16f70363_a0078793,
        64'h67910007_871b0ee6,
        64'h8d63d007_07136725,
        64'h0007869b_0ae68963,
        64'h60070713_67210007,
        64'h869b02d7_68637007,
        64'h07136725_0007869b,
        64'h14e68063_70070713,
        64'h67250007_869baa49,
        64'h14f70863_80078793,
        64'h67890007_871b18e6,
        64'h8b634007_0713670d,
        64'h0007869b_16e68663,
        64'h90070713_67090007,
        64'h869baa7d_16f70763,
        64'h20078793_67850007,
        64'h871b16e6_8e635007,
        64'h07136705_0007869b,
        64'h18e68563_30070713,
        64'h67050007_869b02d7,
        64'h68637007_07136705,
        64'h0007869b_1ae68a63,
        64'h70070713_67050007,
        64'h869b06d7_6c637007,
        64'h0713670d_0007869b,
        64'h20e68463_70070713,
        64'h670d0007_869ba40d,
        64'h1cf70263_b0078793,
        64'h67850007_871b1ce6,
        64'h89636705_0007869b,
        64'h1ce68e63_c0070713,
        64'h67050007_869ba4a9,
        64'h1af70263_70000793,
        64'h0007871b_1ee68563,
        64'h90070713_67050007,
        64'h869b1c07_06632701,
        64'h8007871b_02d76563,
        64'ha0070713_67050007,
        64'h869b20e6_8f63a007,
        64'h07136705_0007869b,
        64'ha47118f7_08633000,
        64'h07930007_871b1ae6,
        64'h85635000_07130007,
        64'h869b2ae6_8e634000,
        64'h07130007_869bac4d,
        64'h18f70d63_10000793,
        64'h0007871b_2c070963,
        64'h0007871b_00d76d63,
        64'h20000713_0007869b,
        64'h1ce68463_20000713,
        64'h0007869b_04d76c63,
        64'h60000713_0007869b,
        64'h20e68563_60000713,
        64'h0007869b_0cd76d63,
        64'h10070713_67050007,
        64'h869b2ae6_8a631007,
        64'h07136705_0007869b,
        64'hfd442783_fef42623,
        64'hfd442783_fcf42a23,
        64'h87aefca4_3c231800,
        64'hf4227179_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623e86f,
        64'he0ef853e_03000593,
        64'h460543dc_fd843783,
        64'hd3a92781_8b85fe04,
        64'h2783a00d_ea4fe0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783fef4_26234789,
        64'he7812781_9bf9fec4,
        64'h2783fef4_262387aa,
        64'he96fe0ef_853e0320,
        64'h059343dc_fd843783,
        64'hc3a12781_8ff967a1,
        64'hfe042703_a899eeef,
        64'he0ef853e_03000593,
        64'h02000613_43dcfd84,
        64'h3783cf81_27810207,
        64'hf7932781_87aaed4f,
        64'he0ef853e_03000593,
        64'h43dcfd84_378302f7,
        64'h1b633007_87936785,
        64'h0007871b_fd442783,
        64'h00f70b63_50078793,
        64'h67850007_871bfd44,
        64'h2783fef4_202387aa,
        64'hf0efe0ef_853e0300,
        64'h059343dc_fd843783,
        64'hef4fe0ef_853a85be,
        64'h27818fd5_2781c467,
        64'hd7831ffe_d7970007,
        64'h869b0107_979bfe44,
        64'h27839301_02079713,
        64'h278127b1_43dcfd84,
        64'h3783a229_fef42623,
        64'h4785c789_27810207,
        64'hf793fe44_2783cb99,
        64'h27818b89_fe842783,
        64'hfef42423_87aaed8f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_02f70f63,
        64'h30078793_67850007,
        64'h871bfd44_278304f7,
        64'h08635007_87936785,
        64'h0007871b_fd442783,
        64'hfef42223_8ff917fd,
        64'h6791fe44_2703fef4,
        64'h222387aa_18c000ef,
        64'hfd843503_85befd44,
        64'h278380bf_e0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'h821fe0ef_853a0300,
        64'h0593fff7_861367c1,
        64'h43d8fd84_3783fd2f,
        64'he0ef853e_85bafd04,
        64'h27039381_17822781,
        64'h27a143dc_fd843783,
        64'h8d1fe0ef_853e02e0,
        64'h05934639_43dcfd84,
        64'h3783863f_e0ef853e,
        64'h4599863a_93411742,
        64'hfcc42703_43dcfd84,
        64'h3783aaed_fef42623,
        64'h4785a419_4785d6e7,
        64'ha2234705_1ffed797,
        64'hca6fe0ef_bb450513,
        64'h00003517_bb458593,
        64'h00003597_44c00613,
        64'ha025cb8d_27818b85,
        64'hfe842783_fef42423,
        64'h87aafe4f_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'hda07a623_1ffed797,
        64'hacb14785_dae7ad23,
        64'h47051ffe_d797cfcf,
        64'he0efc0a5_05130000,
        64'h3517c0a5_85930000,
        64'h359744b0_0613a025,
        64'h04f71e63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_de07a823,
        64'h1ffed797_c385fd84,
        64'h3783fcf4_262387ba,
        64'hfcf42823_87b2fcf4,
        64'h2a238736_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_61457402,
        64'h70a2853e_fec42783,
        64'h0001fcf7_19e301f0,
        64'h07b7873e_27818ff9,
        64'h01f007b7_fe842703,
        64'hfef42423_87aa899f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_a839fef4,
        64'h242387aa_8b7fe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783fcaf_e0ef3e80,
        64'h05139abf_e0ef853a,
        64'h02c00593_863e93c1,
        64'h17c20047_e79393c1,
        64'h17c2fe44_278343d8,
        64'hfd843783_fef42223,
        64'h87aa999f_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783d3ed_27818b89,
        64'hfe442783_fef42223,
        64'h87aa9b9f_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783a821_fef42223,
        64'h87aa9d1f_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783a1bf_e0ef853a,
        64'h02c00593_863e93c1,
        64'h17c20017_e79393c1,
        64'h17c2fe44_278343d8,
        64'hfd843783_fef42223,
        64'h87aaa09f_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783a211_fef42623,
        64'h4785e789_27818ba1,
        64'h2781fe24_5783fef4,
        64'h112387aa_a33fe0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_8a5fe0ef,
        64'h38878513_6785a87f,
        64'he0ef853e_03e00593,
        64'h863afe24_570343dc,
        64'hfd843783_fef41123,
        64'h0087e793_fe245783,
        64'hfef41123_87aaa75f,
        64'he0ef853e_03e00593,
        64'h43dcfd84_3783abff,
        64'he0ef853e_02c00593,
        64'h863afe24_570343dc,
        64'hfd843783_fef41123,
        64'h9be9fe24_5783fef4,
        64'h112387aa_aabfe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_ffe12781,
        64'h8ff901f0_07b7fe84,
        64'h2703fef4_242387aa,
        64'ha33fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783a839,
        64'hfef42423_87aaa51f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_fef42623,
        64'h4785c781_2781fec4,
        64'h2783fef4_262387aa,
        64'h212000ef_fd843503,
        64'hb0078593_67854601,
        64'h4681fca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'hf3e52781_8b892781,
        64'hfeb44783_fef405a3,
        64'h87aabd9f_e0ef853e,
        64'h02f00593_43dcfd84,
        64'h3783a821_fef405a3,
        64'h87aabf1f_e0ef853e,
        64'h02f00593_43dcfd84,
        64'h3783c3bf_e0ef853e,
        64'h02f00593_460943dc,
        64'hfd843783_bcdfe0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783be3f_e0ef853a,
        64'h03000593_fff78613,
        64'h67c143d8_fd843783,
        64'h02e78a23_4709fd84,
        64'h3783a031_02e78a23,
        64'h4705fd84_3783c799,
        64'h2781fec4_2783fef4,
        64'h262387aa_2de000ef,
        64'hfd843503_10000593,
        64'h40ff8637_4681a855,
        64'hfef42623_4785a0c1,
        64'h478510e7_ac234705,
        64'h1ffed797_85bfe0ef,
        64'hf6850513_00003517,
        64'hf6858593_00003597,
        64'h3ac00613_a025cb8d,
        64'h2781fec4_2783fef4,
        64'h262387aa_32e000ef,
        64'hfd843503_45814601,
        64'h4681aa3f_e0ef7107,
        64'h85136789_1607a023,
        64'h1ffed797_aa194785,
        64'h16e7a723_47051ffe,
        64'hd7978b1f_e0effbe5,
        64'h05130000_3517fbe5,
        64'h85930000_35973ab0,
        64'h0613a025_04f71e63,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'h1a07a223_1ffed797,
        64'hc385fd84_3783fca4,
        64'h3c231800_f022f406,
        64'h71798082_614d64ea,
        64'h740a70aa_853efdc4,
        64'h27830001_a0110001,
        64'ha0210001_a031fcf4,
        64'h2e234785_cb892781,
        64'hfdc42783_fcf42e23,
        64'h87aa5100_10eff584,
        64'h35032000_059302f7,
        64'h17634785_873e0347,
        64'hc783f584_378300f7,
        64'h1a634791_873e57fc,
        64'hf5843783_0001a0b9,
        64'hfcf42e23_4785c791,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_7ba020ef,
        64'hf5843503_85befd44,
        64'h2783fcf4_2a231007,
        64'h879b03a2_07b7eb95,
        64'h0a27c783_04c78793,
        64'h1ffed797_a071fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa0ad0_10eff584,
        64'h350302f7_11634791,
        64'h873e57fc_f5843783,
        64'ha865fcf4_2e234785,
        64'h00f70663_4785873e,
        64'h0b97c783_09478793,
        64'h1ffed797_04f71663,
        64'h4791873e_57fcf584,
        64'h378300f7_09634795,
        64'h873e57fc_f5843783,
        64'ha8c5fcf4_2e234785,
        64'h00f70663_4789873e,
        64'h0b97c783_0cc78793,
        64'h1ffed797_02f71063,
        64'h479d873e_57fcf584,
        64'h3783aa29_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h6c4020ef_f5843503,
        64'h10058593_1ffed597,
        64'ha281fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa66b0,
        64'h10eff584_35030cf7,
        64'h0b634799_873e57fc,
        64'hf5843783_d7f84719,
        64'hf5843783_a029d7f8,
        64'h4715f584_378300e7,
        64'hf7634785_873e0377,
        64'hc783f584_3783cf91,
        64'h27818b89_27810c47,
        64'hc7831627_87931ffe,
        64'hd797a825_d7f84711,
        64'hf5843783_00e7f763,
        64'h4785873e_0377c783,
        64'hf5843783_cf912781,
        64'h8bb12781_0c47c783,
        64'h19078793_1ffed797,
        64'ha09dd7f8_471df584,
        64'h378300e7_f7634785,
        64'h873e0377_c783f584,
        64'h3783cf91_27810307,
        64'hf7932781_0c47c783,
        64'h1c078793_1ffed797,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810d47,
        64'hc7831da7_87931ffe,
        64'hd79753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810087,
        64'h979b2781_0d57c783,
        64'h20078793_1ffed797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h8fd92781_0107979b,
        64'h27810d67_c7832267,
        64'h87931ffe_d79753f8,
        64'hf5843783_d3f8f584,
        64'h37830007_871b0187,
        64'h979b2781_0d77c783,
        64'h24878793_1ffed797,
        64'ha461fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa0330,
        64'h20eff584_350326e5,
        64'h85931ffe_d597a47d,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_2cf010ef,
        64'hf5843503_28f71263,
        64'h4795873e_0347c783,
        64'hf5843783_acf1fcf4,
        64'h2e234785_28f70d63,
        64'h4785873e_0b97c783,
        64'h2b878793_1ffed797,
        64'hace5fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa0a30,
        64'h20eff584_35032de5,
        64'h85931ffe_d597ae39,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_048020ef,
        64'hf5843503_d7f84715,
        64'hf5843783_2ee7fd63,
        64'h4785873e_0377c783,
        64'hf5843783_30078563,
        64'h27818b89_27810c47,
        64'hc78332a7_87931ffe,
        64'hd797d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0d47c783_34478793,
        64'h1ffed797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0087979b_27810d57,
        64'hc78336a7_87931ffe,
        64'hd79753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810107,
        64'h979b2781_0d67c783,
        64'h39078793_1ffed797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h0187979b_27810d77,
        64'hc7833b27_87931ffe,
        64'hd797aecd_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h19d020ef_f5843503,
        64'h3d858593_1ffed597,
        64'ha921fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa4390,
        64'h10eff584_350314f7,
        64'h1f634785_873e0367,
        64'hc783f584_378316e7,
        64'hf763478d_873e0357,
        64'hc783f584_378316f7,
        64'h1f634789_873e0347,
        64'hc783f584_3783a19d,
        64'hfcf42e23_47854207,
        64'h83632781_fdc42783,
        64'hfcf42e23_87aa1920,
        64'h20eff584_3503d7f8,
        64'h4715f584_378344e7,
        64'hf3634785_873e0377,
        64'hc783f584_37834407,
        64'h8b632781_8b892781,
        64'hf9d44783_46078263,
        64'h0004c783_02e78e23,
        64'h4705f584_3783fd7f,
        64'he0ef3e80_05139b6f,
        64'hf0ef853a_02c00593,
        64'h863e93c1_17c20047,
        64'he793fda4_578343d8,
        64'hf5843783_fcf41d23,
        64'h87aa9a0f_f0ef853e,
        64'h02c00593_43dcf584,
        64'h3783d3e5_27818b89,
        64'h2781fda4_5783fcf4,
        64'h1d2387aa_9c2ff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_a821fcf4,
        64'h1d2387aa_9daff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_a24ff0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0017e793,
        64'hfda45783_43d8f584,
        64'h3783fcf4_1d2387aa,
        64'ha0eff0ef_853e02c0,
        64'h059343dc_f5843783,
        64'ha3a5fcf4_2e234785,
        64'he7892781_8ba12781,
        64'hfd245783_fcf41923,
        64'h87aaa38f_f0ef853e,
        64'h03e00593_43dcf584,
        64'h37838aaf_f0ef3887,
        64'h85136785_a8cff0ef,
        64'h853e03e0_0593863a,
        64'hfd245703_43dcf584,
        64'h3783fcf4_19230087,
        64'he793fd24_5783fcf4,
        64'h192387aa_a7aff0ef,
        64'h853e03e0_059343dc,
        64'hf5843783_ac4ff0ef,
        64'h853e02c0_0593863a,
        64'hfd245703_43dcf584,
        64'h3783fcf4_19239be9,
        64'hfd245783_fcf41923,
        64'h87aaab0f_f0ef853e,
        64'h02c00593_43dcf584,
        64'h37831407_9d6303c7,
        64'hc783f584_378316f7,
        64'h136347a1_873e4bdc,
        64'hf5843783_16e7fa63,
        64'h478d873e_f9d44783,
        64'h1807d063_4187d79b,
        64'h0187979b_0024c783,
        64'h62079e63_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h19e020ef_f5843503,
        64'h85bef904_0793adb9,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_67f010ef,
        64'hf5843503_c3852781,
        64'h8b912781_0014c783,
        64'ha561fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa4bf0,
        64'h10eff584_350385a6,
        64'ha565fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa3650,
        64'h20eff584_350326f7,
        64'h12634785_873e0347,
        64'hc783f584_3783add9,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_474010ef,
        64'hf5843503_add5fcf4,
        64'h2e234785_adf5fcf4,
        64'h2e234785_cb892781,
        64'hfdc42783_fcf42e23,
        64'h87aa0870_20eff584,
        64'h350385be_5f9cf584,
        64'h3783df98_a807071b,
        64'h018cc737_f5843783,
        64'haf05fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa6e80,
        64'h10eff584_350304f7,
        64'h1b634795_873e0347,
        64'hc783f584_378300f7,
        64'h0a634789_873e0347,
        64'hc783f584_3783a7bd,
        64'hfcf42e23_4785c3d1,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_0f9020ef,
        64'hf5843503_85be5f9c,
        64'hf5843783_df988407,
        64'h071b017d_8737f584,
        64'h3783a801_df98ac07,
        64'h071b0121_f737f584,
        64'h378300f7_1a634789,
        64'h873e0367_c783f584,
        64'h37837c40_006ffcf4,
        64'h2e234785_c7912781,
        64'hfdc42783_fcf42e23,
        64'h87aa915f_f0eff584,
        64'h350306f7_1c634785,
        64'h873e0347_c783f584,
        64'h37837f40_006ffcf4,
        64'h2e234785_00f70763,
        64'h4795873e_0347c783,
        64'hf5843783_00f70f63,
        64'h4789873e_0347c783,
        64'hf5843783_02f70763,
        64'h4785873e_0347c783,
        64'hf5843783_02f702e3,
        64'h47850007_871bfdc4,
        64'h2783fcf4_2e2387aa,
        64'h053000ef_f5843503,
        64'ha83902e7_8a234715,
        64'hf5843783_00f71863,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cf584_37830750,
        64'h006f4785_a4e7a123,
        64'h47051ffe_e797984f,
        64'hf0ef8925_05130000,
        64'h45178925_85930000,
        64'h45972400_0613a02d,
        64'h04f71a63_4789873e,
        64'h0367c783_f5843783,
        64'hdf98a807_071b0006,
        64'h2737f584_37830207,
        64'h8e23f584_378302e7,
        64'h8a234705_f5843783,
        64'h02e78ba3_4705f584,
        64'h3783a807_af231ffe,
        64'he7970e10_006f4785,
        64'haae7a723_47051ffe,
        64'he7979f0f_f0ef8fe5,
        64'h05130000_45178fe5,
        64'h85930000_459723f0,
        64'h0613a02d_06f71963,
        64'h11178793_111117b7,
        64'h873e53dc_f5843783,
        64'hae07a223_1ffee797,
        64'hc385f584_3783fc04,
        64'h3423fc04_3023fa04,
        64'h3c23fa04_3823fa04,
        64'h3423fa04_3023f804,
        64'h3c23f804_38230004,
        64'hb0230057_94938395,
        64'h07fdf807_8793fe04,
        64'h0793f4a4_3c231900,
        64'hed26f122_f5067171,
        64'h80826161_640660a6,
        64'h853efec4_2783fe04,
        64'h2623d3f8_fb843783,
        64'h0007871b_00a7979b,
        64'h27812785_27818ff9,
        64'h17fd0040_07b7873e,
        64'h27810087_d79bfc44,
        64'h278302f7_16634785,
        64'h873e2781_8b8d2781,
        64'h0167d79b_fcc42783,
        64'ha081d3f8_fb843783,
        64'h0007871b_0097d79b,
        64'hfd042783_fcf42823,
        64'h02f707bb_fd842783,
        64'hfd042703_fcf42823,
        64'h02f707bb_fd442703,
        64'h27812785_fd042783,
        64'hfcf42823_8fd9fd04,
        64'h27830007_871b8ff9,
        64'hc0078793_6785873e,
        64'h278100a7_979bfc84,
        64'h2783fcf4_28230167,
        64'hd79bfc44_2783fcf4,
        64'h2a232781_00f717bb,
        64'h47052781_27892781,
        64'h8b9d2781_0077d79b,
        64'hfc442783_fcf42c23,
        64'h278100f7_17bb4705,
        64'h27818bbd_27810087,
        64'hd79bfc84_2783e3c5,
        64'h27818b8d_27810167,
        64'hd79bfcc4_2783fcf4,
        64'h26232781_87aae88f,
        64'hf0ef853e_93811782,
        64'h278127f1_43dcfb84,
        64'h3783fcf4_24232781,
        64'h87aaea4f_f0ef853e,
        64'h93811782_278127e1,
        64'h43dcfb84_3783fcf4,
        64'h22232781_87aaec0f,
        64'hf0ef853e_93811782,
        64'h278127d1_43dcfb84,
        64'h3783fcf4_20232781,
        64'h87aaedcf_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783a28d,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_69f000ef,
        64'hfb843503_90078593,
        64'h6785863e_46814bbc,
        64'hfb843783_d7d54bbc,
        64'hfb843783_cbb8fb84,
        64'h37830007_871b8ff9,
        64'h77c1873e_278187aa,
        64'hf3aff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_a2c1fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa6fd0_00effb84,
        64'h35033000_05934601,
        64'h4681c7f8_fb843783,
        64'h0007871b_87aa81df,
        64'hf0ef853e_45f143dc,
        64'hfb843783_c7b8fb84,
        64'h37830007_871b87aa,
        64'h837ff0ef_853e45e1,
        64'h43dcfb84_3783c3f8,
        64'hfb843783_0007871b,
        64'h87aa851f_f0ef853e,
        64'h45d143dc_fb843783,
        64'hc3b8fb84_37830007,
        64'h871b87aa_86bff0ef,
        64'h853e45c1_43dcfb84,
        64'h3783a4b9_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h78b000ef_fb843503,
        64'h20000593_46014681,
        64'hac95fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa5850,
        64'h00effb84_350302e7,
        64'h8e234705_fb843783,
        64'hc78d2781_8ff90100,
        64'h07b7fe84_2703db98,
        64'h4705fb84_3783c789,
        64'h27818ff9_400007b7,
        64'hfe842703_f407dde3,
        64'hfe842783_fef42423,
        64'h87aa85df_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783a4cd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_01e010ef,
        64'hfb843503_90078593,
        64'h67ad863e_4681fe44,
        64'h2783fef4_22238fd9,
        64'h010007b7_fe442703,
        64'h00f71963_47a1873e,
        64'h4bdcfb84_378302f7,
        64'h10634789_873e0367,
        64'hc783fb84_3783fef4,
        64'h222340ff_87b7a689,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_07e010ef,
        64'hfb843503_70078593,
        64'h678d4601_4681a055,
        64'hfe042423_02e78aa3,
        64'h4709fb84_3783a031,
        64'h02e78aa3_4705fb84,
        64'h378300f7_08631aa0,
        64'h07930007_871bfe84,
        64'h2783fef4_242387aa,
        64'h92bff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_f3e52781,
        64'h8b892781_fe344783,
        64'hfef401a3_87aaa6df,
        64'hf0ef853e_02f00593,
        64'h43dcfb84_3783a821,
        64'hfef401a3_87aaa85f,
        64'hf0ef853e_02f00593,
        64'h43dcfb84_3783acff,
        64'hf0ef853e_02f00593,
        64'h460943dc_fb843783,
        64'h04f71863_47890007,
        64'h871bfec4_2783a129,
        64'hfef42623_478500f7,
        64'h06634789_0007871b,
        64'hfec42783_cf812781,
        64'hfec42783_fef42623,
        64'h87aa1540_10effb84,
        64'h35038007_85936785,
        64'h1aa00613_4681a189,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_17e010ef,
        64'hfb843503_45814601,
        64'h4681a19d_fef42623,
        64'h4785e789_27818ff9,
        64'h67c1fdc4_2703fcf4,
        64'h2e2387aa_a0fff0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfb84,
        64'h3783cb8d_47dcfb84,
        64'h378302f7_0e634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfb843783_a9754785,
        64'hfee7af23_47051ffe,
        64'he797f40f_f0efe4e5,
        64'h05130000_4517e4e5,
        64'h85930000_45971620,
        64'h0613a025_04f71363,
        64'h4789873e_0367c783,
        64'hfb843783_cbd84711,
        64'hfb843783_0207ac23,
        64'h1ffee797_a3114785,
        64'h04e7a323_47051ffe,
        64'he797f88f_f0efe965,
        64'h05130000_4517e965,
        64'h85930000_45971610,
        64'h0613a025_04f71763,
        64'h11178793_111117b7,
        64'h873e53dc_fb843783,
        64'h0607ae23_1ffee797,
        64'hc385fb84_3783faa4,
        64'h3c230880_e0a2e486,
        64'h715d8082_61217442,
        64'h70e2853e_fec42783,
        64'hfe042623_bcdff0ef,
        64'h853e4591_20000613,
        64'h43dcfd84_37830ce7,
        64'h9023474d_1ffee797,
        64'hbe9ff0ef_853e03a0,
        64'h05934601_43dcfd84,
        64'h3783bfbf_f0ef853e,
        64'h03800593_460143dc,
        64'hfd843783_c0dff0ef,
        64'h853a0360_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c23f_f0ef853a,
        64'h03400593_eff78613,
        64'h67c143d8_fd843783,
        64'hcb9ff0ef_853e0280,
        64'h05934641_43dcfd84,
        64'h3783ccbf_f0ef853a,
        64'h02900593_863e0ff7,
        64'hf7930017_e793feb4,
        64'h478343d8_fd843783,
        64'hfe0405a3_a019fef4,
        64'h05a347a9_c7892781,
        64'h8ff90400_07b7873e,
        64'h579cfd84_3783a005,
        64'hfef405a3_47b1c789,
        64'h27818ff9_020007b7,
        64'h873e579c_fd843783,
        64'ha82dfef4_05a347b9,
        64'hc7892781_8ff90100,
        64'h07b7873e_579cfd84,
        64'h3783a8d5_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h154030ef_fd843503,
        64'ha8078593_000627b7,
        64'hb09ff0ef_0c800513,
        64'h00f71663_400007b7,
        64'h873e2781_8ff9c000,
        64'h07b7873e_579cfd84,
        64'h378302f7_13634789,
        64'h873e0367_c783fd84,
        64'h3783d93f_f0ef853e,
        64'h02900593_463d43dc,
        64'hfd843783_a811da7f,
        64'hf0ef853e_02900593,
        64'h463d43dc_fd843783,
        64'h00f71c63_4789873e,
        64'h0367c783_fd843783,
        64'hd798fd84_37830007,
        64'h871b87aa_c7fff0ef,
        64'h853e9381_17822781,
        64'h0407879b_43dcfd84,
        64'h378302e7_8b23fd84,
        64'h37830ff7_f71387aa,
        64'hd3fff0ef_853e0fe0,
        64'h059343dc_fd843783,
        64'hf3e52781_8b852781,
        64'hfea44783_fef40523,
        64'h87aade1f_f0ef853e,
        64'h02f00593_43dcfd84,
        64'h3783a821_fef40523,
        64'h87aadf9f_f0ef853e,
        64'h02f00593_43dcfd84,
        64'h3783e43f_f0ef853e,
        64'h02f00593_460543dc,
        64'hfd843783_bfdff0ef,
        64'h3e800513_e5dff0ef,
        64'h853e0290_05934601,
        64'h43dcfd84_3783a811,
        64'he71ff0ef_853e0290,
        64'h05934641_43dcfd84,
        64'h3783a481_47852ee7,
        64'ha2234705_1ffee797,
        64'ha27ff0ef_13450513,
        64'h00004517_13458593,
        64'h00004597_0b500613,
        64'ha02504f7_10634789,
        64'h873e2781_0ff7f793,
        64'h278187aa_e03ff0ef,
        64'h853e0fe0_059343dc,
        64'hfd843783_0607b823,
        64'hfd843783_d7f84719,
        64'hfd843783_0607a223,
        64'hfd843783_02e78023,
        64'hfd843783_0207c703,
        64'hfd043783_cfd8fd84,
        64'h37834fd8_fd043783,
        64'hcf98fd84_37834f98,
        64'hfd043783_cbd8fd84,
        64'h37834bd8_fd043783,
        64'hcb98fd84_37834b98,
        64'hfd043783_c7d8fd84,
        64'h378347d8_fd043783,
        64'hd3d81117_071b1111,
        64'h1737fd84_3783c798,
        64'hfd843783_4798fd04,
        64'h3783c3d8_fcc42703,
        64'hfd843783_00e79023,
        64'hfd843783_0007d703,
        64'hfd043783_3c07a023,
        64'h1ffee797_a62d4785,
        64'h3ce7a723_47051ffe,
        64'he797b11f_f0ef21e5,
        64'h05130000_451721e5,
        64'h85930000_45970b40,
        64'h0613a025_c7fdfd04,
        64'h37833e07_ab231ffe,
        64'he797cb89_fd843783,
        64'hfcf42623_87b2fcb4,
        64'h3823fca4_3c230080,
        64'hf822fc06_71398082,
        64'h61056442_60e20001,
        64'he8dff0ef_853e85ba,
        64'hfea44703_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h052387ba_fef405a3,
        64'h87b6fef4_26238732,
        64'h86ae87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_853e87aa,
        64'he7fff0ef_853e9381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef405a3_87bafef4,
        64'h2623872e_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e20001,
        64'hf39ff0ef_853e85ba,
        64'hfe845703_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h142387ba_fef405a3,
        64'h87b6fef4_26238732,
        64'h86ae87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_853e87aa,
        64'hf1dff0ef_853e9381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef405a3_87bafef4,
        64'h2623872e_87aa1000,
        64'he822ec06_11018082,
        64'h61457422_0001c398,
        64'hfd442703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf42a23_87aefca4,
        64'h3c231800_f4227179,
        64'h80826145_74220001,
        64'h00e79023_fd645703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf41b23,
        64'h87aefca4_3c231800,
        64'hf4227179_80826145,
        64'h74220001_00e78023,
        64'hfd744703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf40ba3_87aefca4,
        64'h3c231800_f4227179,
        64'h80826105_6462853e,
        64'h2781439c_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61056462,
        64'h853e93c1_17c20007,
        64'hd783fe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826105_6462853e,
        64'h0ff7f793_0007c783,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61457422_853efe84,
        64'h3783fae7_f5e34785,
        64'h0007871b_fe442783,
        64'hfef42223_2785fe44,
        64'h2783a829_fef43423,
        64'h97ba09a7_07130000,
        64'h5717078a_97ba078e,
        64'h87bafe44_670302f7,
        64'h10632781_2701fde4,
        64'h57030007_d78397ba,
        64'h0cc68713_078a97ba,
        64'h078e87ba_fe446703,
        64'h00005697_a0b9fe04,
        64'h2223fe04_3423fcf4,
        64'h1f2387aa_1800f422,
        64'h71798082_61457402,
        64'h70a20001_fef768e3,
        64'hfe043783_fe843703,
        64'hfea43423_fbfff0ef,
        64'hfef43023_97bafe84,
        64'h3783873e_078a97ba,
        64'h078a87ba_fd843703,
        64'hfea43423_fdfff0ef,
        64'hfca43c23_1800f022,
        64'hf4067179_80820141,
        64'h6422853e_639c17e1,
        64'h0200c7b7_0800e422,
        64'h11418082_61096406,
        64'h60a6853e_fec42783,
        64'hfef42623_87aab38f,
        64'hf0efc265_0513ffff,
        64'hf51785be_567dfb84,
        64'h3683fd04_0793fe04,
        64'h3703fcf4_3c23fc04,
        64'h3783fcf4_3823fc84,
        64'h3783fef4_3023fd87,
        64'h87930304_07930314,
        64'h34230304_3023ec1c,
        64'he818e414_fac43c23,
        64'hfcb43023_fca43423,
        64'h0880e0a2_e4867119,
        64'h80826145_740270a2,
        64'h853e87aa_b9eff0ef,
        64'hbf650513_fffff517,
        64'hfe843583_fe043603,
        64'hfd843683_fd043703,
        64'hfcd43823_fcc43c23,
        64'hfeb43023_fea43423,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853e87aa_bdeff0ef,
        64'hc9450513_fffff517,
        64'h85be567d_fd843683,
        64'hfd043703_fe840793,
        64'hfcb43823_fca43c23,
        64'h1800f022_f4067179,
        64'h80826165_744270e2,
        64'h853efec4_2783fef4,
        64'h262387aa_c1eff0ef,
        64'hc7650513_fffff517,
        64'hfd843583_fd043603,
        64'hfc843683_873efe04,
        64'h3783fef4_3023fd87,
        64'h87930304_07930314,
        64'h34230304_3023ec1c,
        64'he818e414_fcc43423,
        64'hfcb43823_fca43c23,
        64'h0080f822_fc067159,
        64'h80826125_740270a2,
        64'h853efec4_2783fef4,
        64'h262387aa_c7eff0ef,
        64'hcd650513_fffff517,
        64'hfd843583_567dfd04,
        64'h3683873e_fe043783,
        64'hfef43023_fd078793,
        64'h03040793_03143423,
        64'h03043023_ec1ce818,
        64'he414e010_fcb43823,
        64'hfca43c23_1800f022,
        64'hf406711d_80826109,
        64'h744270e2_853efec4,
        64'h2783fef4_262387aa,
        64'hcdaff0ef_d9050513,
        64'hfffff517_85be567d,
        64'hfc843683_fd840793,
        64'hfe043703_fef43023,
        64'hfc878793_04040793,
        64'h03143c23_03043823,
        64'hf41cf018_ec14e810,
        64'he40cfca4_34230080,
        64'hf822fc06_71198082,
        64'h610d644a_60ea853e,
        64'h2781fd84_37839702,
        64'h4501f904_3583863e,
        64'hf8843683_f9843703,
        64'hfd843783_a01917fd,
        64'hf8843783_00f76663,
        64'hf8843783_fd843703,
        64'hd8079963_0007c783,
        64'hf8043783_0001f8f4,
        64'h30230785_f8043783,
        64'h9702f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_0007c503,
        64'hf8043783_a80df8f4,
        64'h30230785_f8043783,
        64'h97020250_0513f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'ha8b9f8f4_30230785,
        64'hf8043783_fca43c23,
        64'hba2ff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_87364781,
        64'h484188ba_e03efe84,
        64'h2783e43e_fec42783,
        64'hfe442703_86be639c,
        64'hf6e43c23_00878713,
        64'hf7843783_a089fca4,
        64'h3c23cfcf_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_36838736,
        64'h47814841_88bae03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_270386be,
        64'h639cf6e4_3c230087,
        64'h8713f784_3783c3b1,
        64'h0ff7f793_fbb44783,
        64'hfaf40da3_4785fef4,
        64'h26230217_e793fec4,
        64'h2783fef4_242347c1,
        64'ha239f8f4_30230785,
        64'hf8043783_fce7e7e3,
        64'h2701fe84_2703fce4,
        64'h22230017_871bfc44,
        64'h27839702_02000513,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h3783a00d_cf8d2781,
        64'h8b89fec4_2783fbcd,
        64'hfee42223_fff7871b,
        64'hfe442783_d3e12781,
        64'h4007f793_fec42783,
        64'hcf910007_c783fc84,
        64'h37839702_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_37830007,
        64'hc503fce4_34230017,
        64'h8713fc84_3783a03d,
        64'hfce7e7e3_2701fe84,
        64'h2703fce4_22230017,
        64'h871bfc44_27839702,
        64'h02000513_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_3783a00d,
        64'he7a52781_8b89fec4,
        64'h2783fcf4_222387b2,
        64'h00d77363_0006071b,
        64'h0007869b_fe442783,
        64'hfc442603_cf912781,
        64'h4007f793_fec42783,
        64'hfcf42223_87aa8aaf,
        64'hf0effc84_350385be,
        64'h57fda011_fe446783,
        64'hc7812781_fe442783,
        64'hfcf43423_639cf6e4,
        64'h3c230087_8713f784,
        64'h3783a4a1_f8f43023,
        64'h0785f804_3783fce7,
        64'he7e32701_fe842703,
        64'hfce42823_0017871b,
        64'hfd042783_97020200,
        64'h0513f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_a00dcf8d,
        64'h27818b89_fec42783,
        64'h9702f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_0ff7f513,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783fce7,
        64'he7e32701_fe842703,
        64'hfce42823_0017871b,
        64'hfd042783_97020200,
        64'h0513f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_a00def8d,
        64'h27818b89_fec42783,
        64'hfcf42823_4785a631,
        64'hf8f43023_0785f804,
        64'h3783fca4_3c23e50f,
        64'hf0eff984_3503f904,
        64'h3583fd84_3603f884,
        64'h36834781_883688b2,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442603,
        64'hfd446683_fb446703,
        64'hfaf42a23_2781439c,
        64'hf6e43c23_00878713,
        64'hf7843783_a8012781,
        64'h93c117c2_439cf6e4,
        64'h3c230087_8713f784,
        64'h3783cf81_27810807,
        64'hf793fec4_2783a815,
        64'h27810ff7_f793439c,
        64'hf6e43c23_00878713,
        64'hf7843783_cf812781,
        64'h0407f793_fec42783,
        64'ha841fca4_3c23ee0f,
        64'hf0eff984_3503f904,
        64'h3583fd84_3603f884,
        64'h36834781_883688b2,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442603,
        64'hfd446683_6398f6e4,
        64'h3c230087_8713f784,
        64'h3783c3b1_27811007,
        64'hf793fec4_2783a8f9,
        64'hfca43c23_847ff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h47818836_88b2e03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_2603fd44,
        64'h66836398_f6e43c23,
        64'h00878713_f7843783,
        64'hc3b12781_2007f793,
        64'hfec42783_a235fca4,
        64'h3c23f7cf_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_368387b6,
        64'h883288ae_e03efe84,
        64'h2783e43e_fec42783,
        64'hfe442583_fd446603,
        64'h0ff7f693_01f7d79b,
        64'hfb042783_93010207,
        64'h97132781_278140f7,
        64'h07bb8f3d_fb042703,
        64'h41f7d79b_fb042783,
        64'hfaf42823_439cf6e4,
        64'h3c230087_8713f784,
        64'h3783a801_27814107,
        64'hd79b0107_979b439c,
        64'hf6e43c23_00878713,
        64'hf7843783_cf912781,
        64'h0807f793_fec42783,
        64'ha81d2781_0ff7f793,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783cf81,
        64'h27810407_f793fec4,
        64'h2783a2cd_fca43c23,
        64'h833ff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_872e87ba,
        64'h883688b2_e03efe84,
        64'h2783e43e_fec42783,
        64'hfe442603_fd446683,
        64'h0ff7f713_93fdfa84,
        64'h378385be_8f998fb9,
        64'hfa843783_43f7d713,
        64'hfa843783_faf43423,
        64'h639cf6e4_3c230087,
        64'h8713f784_3783c3bd,
        64'h27811007_f793fec4,
        64'h2783ac89_fca43c23,
        64'h9bbff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_872e87ba,
        64'h883688b2_e03efe84,
        64'h2783e43e_fec42783,
        64'hfe442603_fd446683,
        64'h0ff7f713_93fdfa04,
        64'h378385be_8f998fb9,
        64'hfa043783_43f7d713,
        64'hfa043783_faf43023,
        64'h639cf6e4_3c230087,
        64'h8713f784_3783c3bd,
        64'h27812007_f793fec4,
        64'h278318f7_1d630640,
        64'h0793873e_0007c783,
        64'hf8043783_00f70b63,
        64'h06900793_873e0007,
        64'hc783f804_3783fef4,
        64'h26239bf9_fec42783,
        64'hc7912781_4007f793,
        64'hfec42783_fef42623,
        64'h9bcdfec4_278300f7,
        64'h07630640_0793873e,
        64'h0007c783_f8043783,
        64'h02f70063_06900793,
        64'h873e0007_c783f804,
        64'h3783fef4_26230207,
        64'he793fec4_278300f7,
        64'h18630580_0793873e,
        64'h0007c783_f8043783,
        64'hfef42623_9bbdfec4,
        64'h2783fcf4_2a2347a9,
        64'ha809fcf4_2a234789,
        64'h00f71663_06200793,
        64'h873e0007_c783f804,
        64'h3783a035_fcf42a23,
        64'h47a100f7_166306f0,
        64'h0793873e_0007c783,
        64'hf8043783_a099fcf4,
        64'h2a2347c1_00f71663,
        64'h05800793_873e0007,
        64'hc783f804_378300f7,
        64'h0b630780_0793873e,
        64'h0007c783_f8043783,
        64'h878297ba_ccc78793,
        64'h00005797_0007871b,
        64'h439c97ba_cdc78793,
        64'h00005797_00279713,
        64'h93810206_97936ce7,
        64'he3630530_07930006,
        64'h871bfdb7_869b2781,
        64'h0007c783_f8043783,
        64'h0001a011_0001a021,
        64'h0001a031_f8f43023,
        64'h0785f804_3783fef4,
        64'h26231007_e793fec4,
        64'h2783a015_f8f43023,
        64'h0785f804_3783fef4,
        64'h26231007_e793fec4,
        64'h2783a835_f8f43023,
        64'h0785f804_3783fef4,
        64'h26231007_e793fec4,
        64'h2783a889_f8f43023,
        64'h0785f804_3783fef4,
        64'h26230407_e793fec4,
        64'h278306f7_16630680,
        64'h0793873e_0007c783,
        64'hf8043783_f8f43023,
        64'h0785f804_3783fef4,
        64'h26230807_e793fec4,
        64'h2783a079_f8f43023,
        64'h0785f804_3783fef4,
        64'h26232007_e793fec4,
        64'h27830af7_146306c0,
        64'h0793873e_0007c783,
        64'hf8043783_f8f43023,
        64'h0785f804_3783fef4,
        64'h26231007_e793fec4,
        64'h27838782_97bad927,
        64'h87930000_57970007,
        64'h871b439c_97bada27,
        64'h87930000_57970027,
        64'h97139381_02069793,
        64'h0ee7e963_47c90006,
        64'h871bf987_869b2781,
        64'h0007c783_f8043783,
        64'hf8f43023_0785f804,
        64'h3783fef4_22232781,
        64'h47810007_53630007,
        64'h871bfbc4_2783faf4,
        64'h2e23439c_f6e43c23,
        64'h00878713_f7843783,
        64'h02f71a63_02a00793,
        64'h873e0007_c783f804,
        64'h3783a091_fef42223,
        64'h87aaf86f_f0ef853e,
        64'hf8040793_cb9187aa,
        64'hf54ff0ef_853e0007,
        64'hc783f804_3783f8f4,
        64'h30230785_f8043783,
        64'hfef42623_4007e793,
        64'hfec42783_08f71063,
        64'h02e00793_873e0007,
        64'hc783f804_3783fe04,
        64'h2223f8f4_30230785,
        64'hf8043783_fef42423,
        64'hfc042783_a029fef4,
        64'h24232781_40f007bb,
        64'hfc042783_fef42623,
        64'h0027e793_fec42783,
        64'h0207d063_2781fc04,
        64'h2783fcf4_2023439c,
        64'hf6e43c23_00878713,
        64'hf7843783_04f71763,
        64'h02a00793_873e0007,
        64'hc783f804_3783a8b9,
        64'hfef42423_87aa833f,
        64'hf0ef853e_f8040793,
        64'hcb9187aa_801ff0ef,
        64'h853e0007_c783f804,
        64'h3783fe04_2423f385,
        64'h2781fe04_27830001,
        64'hfe042023_a021fef4,
        64'h20234785_f8f43023,
        64'h0785f804_3783fef4,
        64'h26230107_e793fec4,
        64'h2783a01d_fef42023,
        64'h4785f8f4_30230785,
        64'hf8043783_fef42623,
        64'h0087e793_fec42783,
        64'ha091fef4_20234785,
        64'hf8f43023_0785f804,
        64'h3783fef4_26230047,
        64'he793fec4_2783a08d,
        64'hfef42023_4785f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0027e793,
        64'hfec42783_a041fef4,
        64'h20234785_f8f43023,
        64'h0785f804_3783fef4,
        64'h26230017_e793fec4,
        64'h27838782_97baf467,
        64'h87930000_57970007,
        64'h871b439c_97baf567,
        64'h87930000_57970027,
        64'h97139381_02069793,
        64'h0ce7e063_47c10006,
        64'h871bfe07_869b2781,
        64'h0007c783_f8043783,
        64'hfe042623_f8f43023,
        64'h0785f804_37832270,
        64'h006ff8f4_30230785,
        64'hf8043783_9702f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'h0007c503_f8043783,
        64'h02f70b63_02500793,
        64'h873e0007_c783f804,
        64'h378326b0_006ff8f4,
        64'h3c238667_87930000,
        64'h07972607_9de3f904,
        64'h3783fc04_3c23f6e4,
        64'h3c23f8d4_3023f8c4,
        64'h3423f8b4_3823f8a4,
        64'h3c231100_e922ed06,
        64'h71358082_610d644a,
        64'h60ea853e_87aab47f,
        64'hf0effb84_3503fb04,
        64'h3583fa84_3603fa04,
        64'h3683fe84_37838836,
        64'h88b2e03e_f9042783,
        64'he43e401c_e83e441c,
        64'hfc040713_f9744683,
        64'h0007861b_f8843783,
        64'hf6e7ffe3_47fdfe84,
        64'h3703c791_f9843783,
        64'hf8f43c23_02f757b3,
        64'hf8843783_f9843703,
        64'hfcf70823_9736ff04,
        64'h0693fed4_34230017,
        64'h0693fe84_37030ff7,
        64'hf79337d9_0ff7f793,
        64'h9fb9fe74_47030610,
        64'h0793a019_04100793,
        64'hc7812781_0207f793,
        64'h441ca01d_0ff7f793,
        64'h0307879b_fe744783,
        64'h00e7e963_47a50ff7,
        64'hf713fe74_4783fef4,
        64'h03a302f7_77b3f884,
        64'h3783f984_3703c7c1,
        64'hf9843783_c7812781,
        64'h4007f793_441cc41c,
        64'h9bbd441c_e781f984,
        64'h3783fe04_3423f8f4,
        64'h282387ba_f8f40ba3,
        64'h8746f904_3423f8e4,
        64'h3c23fad4_3023fac4,
        64'h3423fab4_3823faa4,
        64'h3c231100_e922ed06,
        64'h71358082_610d644a,
        64'h60ea853e_87aac5ff,
        64'hf0effb84_3503fb04,
        64'h3583fa84_3603fa04,
        64'h3683fe84_37838836,
        64'h88b2e03e_f9042783,
        64'he43e401c_e83e441c,
        64'hfc040713_f9744683,
        64'h0007861b_f8843783,
        64'hf6e7ffe3_47fdfe84,
        64'h3703c791_f9843783,
        64'hf8f43c23_02f757b3,
        64'hf8843783_f9843703,
        64'hfcf70823_9736ff04,
        64'h0693fed4_34230017,
        64'h0693fe84_37030ff7,
        64'hf79337d9_0ff7f793,
        64'h9fb9fe74_47030610,
        64'h0793a019_04100793,
        64'hc7812781_0207f793,
        64'h441ca01d_0ff7f793,
        64'h0307879b_fe744783,
        64'h00e7e963_47a50ff7,
        64'hf713fe74_4783fef4,
        64'h03a302f7_77b3f884,
        64'h3783f984_3703c7c1,
        64'hf9843783_c7812781,
        64'h4007f793_441cc41c,
        64'h9bbd441c_e781f984,
        64'h3783fe04_3423f8f4,
        64'h282387ba_f8f40ba3,
        64'h8746f904_3423f8e4,
        64'h3c23fad4_3023fac4,
        64'h3423fab4_3823faa4,
        64'h3c231100_e922ed06,
        64'h71358082_61616406,
        64'h60a6853e_87aac65f,
        64'hf0effe84_3503fe04,
        64'h3583fd84_3603fd04,
        64'h3683fc84_3703fc04,
        64'h3783883e_88ba441c,
        64'h481800e7_80230200,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_cf912781,
        64'h8ba1481c_a01500e7,
        64'h802302b0_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'hcf992781_8b91481c,
        64'ha0a100e7_802302d0,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_cf990ff7,
        64'hf793fbf4_478306e7,
        64'he86347fd_fc043703,
        64'h00e78023_03000713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h378300e7_ef6347fd,
        64'hfc043703_00e78023,
        64'h06200713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_378300e7,
        64'hef6347fd_fc043703,
        64'h02f71463_47890007,
        64'h871bfb84_2783a815,
        64'h00e78023_05800713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h378302e7_e06347fd,
        64'hfc043703_c7852781,
        64'h0207f793_481c02f7,
        64'h1a6347c1_0007871b,
        64'hfb842783_a88d00e7,
        64'h80230780_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'h02e7e063_47fdfc04,
        64'h3703e785_27810207,
        64'hf793481c_02f71a63,
        64'h47c10007_871bfb84,
        64'h2783fcf4_302317fd,
        64'hfc043783_00f71763,
        64'h47c10007_871bfb84,
        64'h2783cf89_fc043783,
        64'hfcf43023_17fdfc04,
        64'h378302f7_1663fc04,
        64'h37030084_678300f7,
        64'h0863fc04_37030004,
        64'h6783c3a9_fc043783,
        64'he7a12781_4007f793,
        64'h481c1207_83632781,
        64'h8bc1481c_fce7f6e3,
        64'h47fdfc04_370300f7,
        64'h7763fc04_37030084,
        64'h6783cf81_27818b85,
        64'h481c00e7_80230300,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_a831fce7,
        64'hfae347fd_fc043703,
        64'h02f77563_fc043703,
        64'h00046783_00e78023,
        64'h03000713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_3783a831,
        64'hc41c37fd_441cc395,
        64'h27818bb1_481ce789,
        64'h0ff7f793_fbf44783,
        64'hcb9d2781_8b85481c,
        64'hcf9d2781_441cebd1,
        64'h27818b89_481cfaf4,
        64'h2c2387ba_faf40fa3,
        64'h874687c2_fcf43023,
        64'hfce43423_fcd43823,
        64'hfcc43c23_feb43023,
        64'hfea43423_0880e0a2,
        64'he486715d_80826125,
        64'h644660e6_853efc84,
        64'h3783fcf7_69e3fac4,
        64'h67838f1d_fe043783,
        64'hfc843703_97020200,
        64'h0513fd04_3583863e,
        64'hfc043683_fd843703,
        64'hfce43423_00178713,
        64'hfc843783_a00dcb9d,
        64'h27818b89_fa842783,
        64'hf7e1fb04_37839702,
        64'hfd043583_863efc04,
        64'h3683fd84_3703fce4,
        64'h34230017_8713fc84,
        64'h37830007_c50397ba,
        64'hfb043783_fb843703,
        64'hfaf43823_17fdfb04,
        64'h3783a81d_fcf767e3,
        64'hfe843703_fac46783,
        64'hfef43423_0785fe84,
        64'h37839702_02000513,
        64'hfd043583_863efc04,
        64'h3683fd84_3703fce4,
        64'h34230017_8713fc84,
        64'h3783a035_fef43423,
        64'hfb043783_efa52781,
        64'h8b85fa84_2783e3c9,
        64'h27818b89_fa842783,
        64'hfef43023_fc843783,
        64'hfaf42423_87bafaf4,
        64'h26238746_87c2faf4,
        64'h3823fae4_3c23fcd4,
        64'h3023fcc4_3423fcb4,
        64'h3823fca4_3c231080,
        64'he8a2ec86_711d8082,
        64'h61457402_70a2853e,
        64'hfec42783_ffc587aa,
        64'hf6dff0ef_853e0007,
        64'hc783639c_fd843783,
        64'hfef42623_fd07879b,
        64'h27819fb9_27810007,
        64'hc783e290_fd843683,
        64'h00178613_639cfd84,
        64'h37830007_871b0017,
        64'h979b9fb9_0027979b,
        64'h87bafec4_2703a825,
        64'hfe042623_fca43c23,
        64'h1800f022_f4067179,
        64'h80826105_6462853e,
        64'h0ff7f793_8b854781,
        64'ha0114785_00e7e463,
        64'h03900793_0ff7f713,
        64'hfef44783_00e7fc63,
        64'h02f00793_0ff7f713,
        64'hfef44783_fef407a3,
        64'h87aa1000_ec221101,
        64'h80826145_7422853e,
        64'h278140f7_07b3fd84,
        64'h3783fe84_3703f3e5,
        64'hfce43823_fff78713,
        64'hfd043783_cb810007,
        64'hc783fe84_3783fef4,
        64'h34230785_fe843783,
        64'ha031fef4_3423fd84,
        64'h3783fcb4_3823fca4,
        64'h3c231800_f4227179,
        64'h80826145_740270a2,
        64'h00019682_853e85ba,
        64'hfef44783_6798fe04,
        64'h37836394_fe043783,
        64'hcf810ff7_f793fef4,
        64'h4783fef4_07a3fcd4,
        64'h3823fcc4_3c23feb4,
        64'h302387aa_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_0001959f,
        64'hf0ef853e_fef44783,
        64'hc7910ff7_f793fef4,
        64'h4783fef4_07a3fcd4,
        64'h3823fcc4_3c23feb4,
        64'h302387aa_1800f022,
        64'hf4067179_80826145,
        64'h74220001_fef407a3,
        64'hfcd43823_fcc43c23,
        64'hfeb43023_87aa1800,
        64'hf4227179_80826145,
        64'h74220001_00e78023,
        64'hfef44703_97bafd84,
        64'h3783fe04_370300f7,
        64'h7b63fd04_3783fd84,
        64'h3703fef4_07a3fcd4,
        64'h3823fcc4_3c23feb4,
        64'h302387aa_1800f422,
        64'h71798082_610d690a,
        64'h64aa644a_60eaf604,
        64'h0113853e_8126814a,
        64'h47812b00_10ef7ce5,
        64'h05130000_5517a801,
        64'h57f92c00_10ef58e5,
        64'h05130000_551785be,
        64'hfac42783_2d2010ef,
        64'h58850513_00005517,
        64'hc3952781_fac42783,
        64'hfaf42623_87aabd5f,
        64'hf0eff684_350385be,
        64'h863af644_27032781,
        64'h739cf804_37833040,
        64'h10ef80a5_05130000,
        64'h6517f8f4_3023f884,
        64'h3783eae7_d2e3478d,
        64'h0007871b_fd042783,
        64'hfcf42823_2785fd04,
        64'h27833300_10ef6565,
        64'h05130000_5517fce7,
        64'hd6e30470_07930007,
        64'h871bfdc4_2783fcf4,
        64'h2e232785_fdc42783,
        64'h356010ef_7d450513,
        64'h00005517_85be2781,
        64'h0387c783_97bafdc4,
        64'h2783f784_3703a02d,
        64'hfc042e23_37a010ef,
        64'h86850513_00006517,
        64'h386010ef_85c50513,
        64'h00006517_85be7b9c,
        64'hf7843783_39a010ef,
        64'h85850513_00006517,
        64'h85be779c_f7843783,
        64'h3ae010ef_85450513,
        64'h00006517_85be739c,
        64'hf7843783_fce7d7e3,
        64'h47bd0007_871bfd84,
        64'h2783fcf4_2c232785,
        64'hfd842783_3da010ef,
        64'h85850513_00006517,
        64'h85be2781_0107c783,
        64'h97bafd84_2783f784,
        64'h3703a02d_fc042c23,
        64'h3fe010ef_88450513,
        64'h00006517_fce7d7e3,
        64'h47bd0007_871bfd44,
        64'h2783fcf4_2a232785,
        64'hfd442783_422010ef,
        64'h8a050513_00006517,
        64'h85be2781_0007c783,
        64'h97bafd44_2783f784,
        64'h3703a02d_fc042a23,
        64'h446010ef_8a450513,
        64'h00006517_452010ef,
        64'h89850513_00006517,
        64'h85befd04_2783f6f4,
        64'h3c2397ba_27010077,
        64'h171bfd04_2703f884,
        64'h3783aa91_fc042823,
        64'haac957f9_482010ef,
        64'h8a850513_00006517,
        64'h85befac4_27834940,
        64'h10ef74a5_05130000,
        64'h5517c395_2781fac4,
        64'h2783faf4_262387aa,
        64'hd97ff0ef_853a85be,
        64'h46052781_67bcfa04,
        64'h3783f884_3703f8f4,
        64'h34230007_8793878a,
        64'h40f10133_07928391,
        64'h07bdf8e4_3823177d,
        64'h873e893a_870afc04,
        64'h37834e80_10ef8ee5,
        64'h05130000_651785be,
        64'h4bfcfa04_37834fc0,
        64'h10ef8e25_05130000,
        64'h651785be_4bbcfa04,
        64'h37835100_10ef8ce5,
        64'h05130000_651785be,
        64'h67bcfa04_37835240,
        64'h10ef8ca5_05130000,
        64'h651785be_739cfa04,
        64'h37835380_10ef8c65,
        64'h05130000_651785be,
        64'h6f9cfa04_378354c0,
        64'h10ef8c25_05130000,
        64'h651785be_4bdcfa04,
        64'h37835600_10ef8be5,
        64'h05130000_651785be,
        64'h4b9cfa04_37835740,
        64'h10ef8ba5_05130000,
        64'h651785be_47dcfa04,
        64'h37835880_10ef8b65,
        64'h05130000_651785be,
        64'h479cfa04_378359c0,
        64'h10ef8c25_05130000,
        64'h6517fce7_d7e3479d,
        64'h0007871b_fcc42783,
        64'hfcf42623_2785fcc4,
        64'h27835c00_10ef8de5,
        64'h05130000_651785be,
        64'h27810007_c78397ba,
        64'hf9843703_fcc42783,
        64'ha02dfc04_2623f8f4,
        64'h3c23fa04_37835ec0,
        64'h10ef8fa5_05130000,
        64'h65175f80_10ef8e65,
        64'h05130000_6517faf4,
        64'h3023fb04_3783a68d,
        64'h57f96100_10ef8de5,
        64'h05130000_651785be,
        64'hfac42783_622010ef,
        64'h8d850513_00006517,
        64'hc3952781_fac42783,
        64'hfaf42623_87aaf25f,
        64'hf0ef853e_45854605,
        64'hfb043783_faf43823,
        64'h00078793_878a40f1,
        64'h01330792_839107bd,
        64'hfae43c23_177d873e,
        64'hfc043783_fcf43023,
        64'h20000793_672010ef,
        64'h91050513_00006517,
        64'haed157fd_682010ef,
        64'h8f850513_00006517,
        64'hcb892781_fc842783,
        64'hfcf42423_87aaecdf,
        64'hf0ef84be_878af6f4,
        64'h222387ae_f6a43423,
        64'h1100e14a_e526e922,
        64'hed067135_80826145,
        64'h740270a2_853e4781,
        64'ha01157fd_6ca010ef,
        64'h92050513_00006517,
        64'h85befec4_2783cf81,
        64'h2781fec4_2783fef4,
        64'h262387aa_7b8030ef,
        64'hc3050513_1fff0517,
        64'h85be4605_fd843683,
        64'hfd442783_fcf42823,
        64'h87bafcf4_2a238732,
        64'h87aefca4_3c231800,
        64'hf022f406_71798082,
        64'h61056442_60e2853e,
        64'h47817280_10ef95e5,
        64'h05130000_6517a801,
        64'h57f57380_10ef93e5,
        64'h05130000_651785be,
        64'hfe442783_cf812781,
        64'hfe442783_fef42223,
        64'h87aa4ee0_20efc9e5,
        64'h05131fff_0517a081,
        64'h57f97680_10ef9465,
        64'h05130000_651785be,
        64'hfe442783_cf812781,
        64'hfe442783_fef42223,
        64'h87aa4390_10efcce5,
        64'h05131fff_0517fe84,
        64'h3583863e_43dcfe84,
        64'h3783a8b5_57fd7a40,
        64'h10ef9625_05130000,
        64'h6517eb89_fe843783,
        64'hfea43423_217010ef,
        64'h45017c00_10ef9665,
        64'h05130000_65171000,
        64'he822ec06_11018082,
        64'h61457402_70a20001,
        64'heb9ff0ef_01078513,
        64'h07fa478d_02000593,
        64'hec9ff0ef_00878513,
        64'h07fa478d_0c700593,
        64'hed9ff0ef_00c78513,
        64'h07fa478d_458dee7f,
        64'hf0ef0047_851307fa,
        64'h478d85be_0ff7f793,
        64'h27810087_d79bfec4,
        64'h2783f03f_f0ef01e7,
        64'h9513478d_85be0ff7,
        64'hf793fec4_2783f17f,
        64'hf0ef00c7_851307fa,
        64'h478d0800_0593f27f,
        64'hf0ef0047_851307fa,
        64'h478d4581_fef42623,
        64'h02f757bb_fdc42703,
        64'h27810047_979bfd84,
        64'h2783fcf4_2c2387ba,
        64'hfcf42e23_872e87aa,
        64'h1800f022_f4067179,
        64'h80826105_644260e2,
        64'h0001f6bf_f0ef01e7,
        64'h9513478d_85befef4,
        64'h4783dfed_87aafc9f,
        64'hf0ef0001_fef407a3,
        64'h87aa1000_e822ec06,
        64'h11018082_01416402,
        64'h60a2853e_27810207,
        64'hf7932781_87aafd3f,
        64'hf0ef0147_851307fa,
        64'h478d0800_e022e406,
        64'h11418082_61056462,
        64'h853e0ff7_f7930007,
        64'hc783fe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826145_74220001,
        64'h00e78023_fd744703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf40ba3,
        64'h87aefca4_3c231800,
        64'hf4227179_a00112d0,
        64'h10efaaa5_05130000,
        64'h65178402_07c58593,
        64'h00006597_10000437,
        64'heb812781_fe842783,
        64'hfef42423_87aa29e0,
        64'h00ef1000_053765a1,
        64'h15f010ef_ad450513,
        64'h00006517_fce7dae3,
        64'h47890007_871bfec4,
        64'h2783fef4_26232785,
        64'hfec42783_183010ef,
        64'haf050513_00006517,
        64'h3a1010ef_24078513,
        64'h000f47b7_a015fe04,
        64'h26231a10_10efae65,
        64'h05130000_651712a0,
        64'h00efa007_85130262,
        64'h67b72007_859367f1,
        64'h1000e822_ec061101,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00048067,
        64'h100004b7_18458593,
        64'h00006597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h0e4000ef_fec10113,
        64'h3fff0117_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
