/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 3529;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_322d746c,
        64'h75616665_642d6972,
        64'h742c786e_6c780074,
        64'h6c756166_65642d69,
        64'h72742c78_6e6c7800,
        64'h6c617564_2d73692c,
        64'h786e6c78_00746e65,
        64'h73657270_2d747075,
        64'h72726574_6e692c78,
        64'h6e6c7800_68746469,
        64'h772d326f_6970672c,
        64'h786e6c78_00687464,
        64'h69772d6f_6970672c,
        64'h786e6c78_00322d74,
        64'h6c756166_65642d74,
        64'h756f642c_786e6c78,
        64'h00746c75_61666564,
        64'h2d74756f_642c786e,
        64'h6c780032_2d737475,
        64'h706e692d_6c6c612c,
        64'h786e6c78_00737475,
        64'h706e692d_6c6c612c,
        64'h786e6c78_0072656c,
        64'h6c6f7274_6e6f632d,
        64'h6f697067_00736c6c,
        64'h65632d6f_69706723,
        64'h0070772d_656c6261,
        64'h73696400_7365676e,
        64'h61722d65_6761746c,
        64'h6f760079_636e6575,
        64'h71657266_2d78616d,
        64'h2d697073_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_5a020000,
        64'h04000000_03000000,
        64'hffffffff_49020000,
        64'h04000000_03000000,
        64'h01000000_3c020000,
        64'h04000000_03000000,
        64'h00000000_25020000,
        64'h04000000_03000000,
        64'h08000000_14020000,
        64'h04000000_03000000,
        64'h08000000_04020000,
        64'h04000000_03000000,
        64'h00000000_f0010000,
        64'h04000000_03000000,
        64'h00000000_de010000,
        64'h04000000_03000000,
        64'h00000000_cc010000,
        64'h04000000_03000000,
        64'h00000000_bc010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h000000c1_00000000,
        64'h67000000_10000000,
        64'h03000000_ac010000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'ha0010000_04000000,
        64'h03000000_00000030,
        64'h30303030_30316340,
        64'h6f697067_01000000,
        64'h02000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_03000000,
        64'h52010000_04000000,
        64'h03000000_00000000,
        64'h64656c62_61736964,
        64'h6b000000_09000000,
        64'h03000000_00100000,
        64'h00000000_00b000e0,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00006d65_672c736e,
        64'h6463006d_65672d71,
        64'h6e797a2c_736e6463,
        64'h1b000000_17000000,
        64'h03000000_00000030,
        64'h30306230_30306540,
        64'h74656e72_65687465,
        64'h01000000_02000000,
        64'h02000000_95010000,
        64'h00000000_03000000,
        64'he40c0000_e40c0000,
        64'h86010000_08000000,
        64'h03000000_20bcbe00,
        64'h74010000_04000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00000000,
        64'h746f6c73_2d697073,
        64'h2d636d6d_1b000000,
        64'h0d000000_03000000,
        64'h00000030_40636d6d,
        64'h01000000_00100000,
        64'h00000000_000010e0,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_52010000,
        64'h04000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h00000000_64656c62,
        64'h61736964_6b000000,
        64'h09000000_03000000,
        64'h00000061_392e382d,
        64'h69636864_732c6e61,
        64'h73617261_1b000000,
        64'h12000000_03000000,
        64'h00000000_30303030,
        64'h30313065_40636d6d,
        64'h01000000_02000000,
        64'h00100000_00000000,
        64'h00d000e0_00000000,
        64'h67000000_10000000,
        64'h03000000_02000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h64656c62_61736964,
        64'h6b000000_09000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_0000302e,
        64'h312d6970_73712d71,
        64'h6e797a2c_786e6c78,
        64'h1b000000_13000000,
        64'h03000000_00000000,
        64'h30303064_30303065,
        64'h40697073_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_005a6202,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_000000c0,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30306340,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000030_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h31407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_005a6202,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30634074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08090000_6d020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h40090000_38000000,
        64'had0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'hffffb3f2_ffffba8e,
        64'hffffba8e_ffffb3f2,
        64'hffffba8e_ffffb878,
        64'hffffba8e_ffffba8e,
        64'hffffb9b2_ffffb3f2,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffb3f2,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffb3f2_ffffb7b4,
        64'hffffb3f2_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffb3f2_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba8e,
        64'hffffba8e_ffffba62,
        64'hffffb3dc_ffffb3f4,
        64'hffffb3f4_ffffb3f4,
        64'hffffb3f4_ffffb3f4,
        64'hffffb3ac_ffffb3f4,
        64'hffffb3f4_ffffb3f4,
        64'hffffb3f4_ffffb3f4,
        64'hffffb3f4_ffffb3f4,
        64'hffffb32c_ffffb3f4,
        64'hffffb3c4_ffffb3f4,
        64'hffffb36c_ffffb178,
        64'hffffb20e_ffffb20e,
        64'hffffb196_ffffb20e,
        64'hffffb1b4_ffffb20e,
        64'hffffb20e_ffffb20e,
        64'hffffb20e_ffffb20e,
        64'hffffb20e_ffffb20e,
        64'hffffb1f0_ffffb20e,
        64'hffffb20e_ffffb1d2,
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00586c6c_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000000_00007525,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000000_00007525,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_58323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h000a5838_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h000a5838_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_000a586c,
        64'h6c363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h00000000_0a756c6c,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h00000000_0a756c6c,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_0a583830,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_0a583830,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_0a583830,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_0a583830,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h00000000_0000000a,
        64'h00000000_00006325,
        64'h00202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h00000000_0a642520,
        64'h3a737574_61747320,
        64'h2c64656c_69616620,
        64'h64616552_20304453,
        64'h00000000_0a216465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a6425,
        64'h203a7375_74617473,
        64'h202c6465_6c696166,
        64'h206e6f69_74617a69,
        64'h6c616974_696e6920,
        64'h64726163_20304453,
        64'h0000000a_6425203a,
        64'h73757461_7473202c,
        64'h64656c69_6166206c,
        64'h61697469_6e692067,
        64'h69666e6f_63204453,
        64'h00000000_0000000a,
        64'h2164656c_69616620,
        64'h6769666e_6f632070,
        64'h756b6f6f_6c204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000020_58323025,
        64'h00000000_0000000a,
        64'h786c6c25_78304045,
        64'h5341425f_4d415244,
        64'h00000000_0000000a,
        64'h00000000_002e2e2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623a14f_c0ef4505,
        64'ha031fef4_26234785,
        64'he7892781_0807f793,
        64'h278187aa_aa5fe0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_0001a011,
        64'hf6e7fee3_02700793,
        64'h0ff7f713_fe944783,
        64'hfef404a3_2785fe94,
        64'h4783cf99_27810407,
        64'hf7932781_87aaadff,
        64'he0ef853e_03e00593,
        64'h43dcfd84_3783a0ad,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_ae5fd0ef,
        64'hfd843503_50078593,
        64'h67854601_4685a829,
        64'hfef42623_87aaafff,
        64'hd0effd84_35033007,
        64'h85936785_46014685,
        64'h00f71f63_4785873e,
        64'h0347c783_fd843783,
        64'ha8adfe04_04a3ad0f,
        64'hc0ef4505_b87fe0ef,
        64'h853e03e0_0593863a,
        64'hfe645703_43dcfd84,
        64'h3783fef4_13230407,
        64'he793fe64_5783fef4,
        64'h132387aa_b75fe0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_c4e19023,
        64'h4741bc5f_e0ef853e,
        64'h4591863a_fea45703,
        64'h43dcfd84_3783fef4,
        64'h15238ff9_17fd6785,
        64'hfea45703_fef41523,
        64'h0017979b_fea45783,
        64'haa254785_c2e1ae23,
        64'h470593af_c0ef7b65,
        64'h05130000_05177ae5,
        64'h85930000_05974b60,
        64'h0613a015_02f71a63,
        64'h478d873e_0377c783,
        64'hfd843783_fef41523,
        64'h04000793_c201ae23,
        64'haaa54785_c2e1ae23,
        64'h470597af_c0ef7f65,
        64'h05130000_05177ee5,
        64'h85930000_05974b50,
        64'h0613a015_04f71363,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'hc201ae23_cf91fd84,
        64'h3783fca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'hbeffe0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_caffe0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe842783,
        64'ha83dfef4_26234785,
        64'hcd3fe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe84,
        64'h2703fef4_242387aa,
        64'hcc1fe0ef_853e0300,
        64'h059343dc_fd843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aacc7f,
        64'hd0effd84_35036000,
        64'h0593863e_4681fd44,
        64'h2783fcf4_2a2387ae,
        64'hfca43c23_1800f022,
        64'hf4067179_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aacb5f,
        64'he0ef853e_93811782,
        64'h278127c1_43dcfc84,
        64'h3783d75f_e0ef853e,
        64'h03000593_460943dc,
        64'hfc843783_dfc52781,
        64'h8b89fdc4_2783a83d,
        64'hfef42623_4785d99f,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfc843783_c3852781,
        64'h8ff967a1_fdc42703,
        64'hfcf42e23_87aad87f,
        64'he0ef853e_03000593,
        64'h43dcfc84_3783a8bd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_d8dfd0ef,
        64'hfc843503_80078593,
        64'h6785863e_4685fe44,
        64'h2783c4e1_90234745,
        64'h7010d073_70105073,
        64'h0ff0000f_fc2fe0ef,
        64'hfc843503_85befc04,
        64'h36032781_fe245783,
        64'he23fe0ef_853e4591,
        64'h863afe04_570343dc,
        64'hfc843783_fef41023,
        64'h8ff917fd_6785fe04,
        64'h5703fef4_10232000,
        64'h0793fef4_11234785,
        64'hfce7dee3_1ff00793,
        64'h0007871b_fe842783,
        64'hfef42423_2785fe84,
        64'h27830007_802397ba,
        64'hfc043703_fe842783,
        64'ha2354785_c2e1ae23,
        64'h4705bc2f_c0efa3e5,
        64'h05130000_1517a365,
        64'h85930000_15973750,
        64'h0613a835_fe042423,
        64'hc201ae23_aaa14785,
        64'hc2e1ae23_4705beef,
        64'hc0efa6a5_05130000,
        64'h1517a625_85930000,
        64'h15973740_0613a015,
        64'h02f71963_11178793,
        64'h111117b7_873e53dc,
        64'hfc843783_c201ae23,
        64'hcf91fc84_3783fe04,
        64'h2223fcb4_3023fca4,
        64'h34230080_f822fc06,
        64'h71398082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_a019fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaecbf_d0effd84,
        64'h3503a007_859367ad,
        64'h46014681_a03dfef4,
        64'h26234785_a82d4785,
        64'hc2e1ae23_4705c86f,
        64'hc0efb025_05130000,
        64'h1517afa5_85930000,
        64'h15973450_0613a015,
        64'hc79d2781_fec42783,
        64'hfef42623_87aaf17f,
        64'hd0effd84_35037007,
        64'h8593678d_863e4681,
        64'h4bbcfd84_3783c201,
        64'hae23a061_4785c2e1,
        64'hae234705_cd4fc0ef,
        64'hb5050513_00001517,
        64'hb4858593_00001597,
        64'h34400613_a01504f7,
        64'h1a631117_87931111,
        64'h17b7873e_53dcfd84,
        64'h3783c201_ae23cf91,
        64'hfd843783_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efe84_2783fe04,
        64'h2423fedf_e0ef853a,
        64'h02c00593_863e93c1,
        64'h17c20047_e793fe44,
        64'h578343d8_fd843783,
        64'hfef41223_87aafd7f,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783d3e5,
        64'h27818b89_2781fe64,
        64'h5783fef4_132387aa,
        64'hff9fe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'ha821fef4_132387aa,
        64'h810ff0ef_853e02c0,
        64'h059343dc_fd843783,
        64'h85aff0ef_853e02c0,
        64'h0593863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12230017_e79393c1,
        64'h17c28fd9_fe445783,
        64'hfec45703_fef41623,
        64'hf007f793_fec45783,
        64'hfef41623_0087979b,
        64'hfec45783_fef41223,
        64'h0ff7f793_fe445783,
        64'hfef41223_87aa876f,
        64'hf0ef853e_02c00593,
        64'h43dcfd84_3783a0a5,
        64'h8c2ff0ef_853e02c0,
        64'h0593863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12230017_e79393c1,
        64'h17c28fd9_fe445783,
        64'h93410307_97138fd9,
        64'hfe245783_fec45703,
        64'hfef41623_f007f793,
        64'hfec45783_fef41623,
        64'h0087979b_fec45783,
        64'hfef41123_0c07f793,
        64'hfe245783_fef41123,
        64'h0067979b_fe245783,
        64'hfef41123_0087d79b,
        64'hfec45783_fef41223,
        64'h03f7f793_fe445783,
        64'hfef41223_87aa90ef,
        64'hf0ef853e_02c00593,
        64'h43dcfd84_378308f7,
        64'h1e634789_873e0367,
        64'hc783fd84_3783a249,
        64'hfef42423_478500e7,
        64'hf6631000_07930007,
        64'h871bfee4_5783fae7,
        64'hfee31000_07930007,
        64'h871bfee4_5783fef4,
        64'h17230017_979bfee4,
        64'h5783a839_fef41623,
        64'h0017d79b_fee45783,
        64'h00e7e963_2781fd44,
        64'h27830007_871b02f7,
        64'h57bb2781_fee45783,
        64'h4798fd84_3783a82d,
        64'hfef41723_4785a2ed,
        64'hfef42423_478506e7,
        64'hfa637fe0_07930007,
        64'h871bfee4_5783fae7,
        64'hffe37fe0_07930007,
        64'h871bfee4_5783fef4,
        64'h17232785_fee45783,
        64'ha831fef4_16230017,
        64'hd79bfee4_578300e7,
        64'he9632781_fd442783,
        64'h0007871b_02f757bb,
        64'h2781fee4_57834798,
        64'hfd843783_a825fef4,
        64'h17234785_ac914785,
        64'hc2e1ae23_4705f7ef,
        64'hc0efdfa5_05130000,
        64'h1517df25_85930000,
        64'h15972d00_0613a015,
        64'h08f71763_4789873e,
        64'h0367c783_fd843783,
        64'ha6aff0ef_853e02c0,
        64'h0593863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12239be9_fe445783,
        64'hfef41223_87aaa56f,
        64'hf0ef853e_02c00593,
        64'h43dcfd84_3783c201,
        64'hae23a4c9_4785c2e1,
        64'hae234705_fecfc0ef,
        64'he6850513_00001517,
        64'he6058593_00001597,
        64'h2cf00613_a01506f7,
        64'h1a631117_87931111,
        64'h17b7873e_53dcfd84,
        64'h3783c201_ae23cf91,
        64'hfd843783_fe041623,
        64'hfcf42a23_87aefca4,
        64'h3c231800_f022f406,
        64'h71798082_61657406,
        64'h70a6853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_a6aff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_f9843783,
        64'hbaaff0ef_853e0280,
        64'h0593863a_0ff77713,
        64'hfe442703_43dcf984,
        64'h3783fef4_22230047,
        64'he793fe44_2783fef4,
        64'h222387aa_b9cff0ef,
        64'h853e0280_059343dc,
        64'hf9843783_ab7fc0ef,
        64'h3e800513_a09dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa7080_00eff984,
        64'h350302f7_1163479d,
        64'h873e57fc_f9843783,
        64'ha849fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa0b80,
        64'h00eff984_350385be,
        64'h5f9cf984_3783bc0f,
        64'hf0ef853e_03000593,
        64'h460943dc_f9843783,
        64'hdfc52781_8b89fe44,
        64'h2783a8d1_fef42623,
        64'h4785be4f_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_f9843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aabd2f_f0ef853e,
        64'h03000593_43dcf984,
        64'h3783aa11_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hbd8fe0ef_f9843503,
        64'h60000593_863e4681,
        64'hfe842783_df985007,
        64'h071b0319_7737f984,
        64'h3783fef4_24231007,
        64'h879b03b9_07b7a831,
        64'hdf985007_071b0319,
        64'h7737f984_3783fef4,
        64'h24231007_879b03b9,
        64'h07b702f7_10634791,
        64'h873e57fc_f9843783,
        64'ha099df98_2007071b,
        64'h0bebc737_f9843783,
        64'hfef42423_2007879b,
        64'h03b907b7_02f71063,
        64'h479d873e_57fcf984,
        64'h3783a275_fef42623,
        64'h47851407_89632781,
        64'hfec42783_fef42623,
        64'h87aa1d40_00eff984,
        64'h35035007_85930319,
        64'h77b7df98_5007071b,
        64'h03197737_f9843783,
        64'hceaff0ef_853e0300,
        64'h05934609_43dcf984,
        64'h3783dfc5_27818b89,
        64'hfe442783_aafdfef4,
        64'h26234785_d0eff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8f984,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_cfcff0ef,
        64'h853e0300_059343dc,
        64'hf9843783_ac3dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aad02f_e0eff984,
        64'h35036000_0593863e,
        64'h4681fe84_2783fef4,
        64'h24231007_879b03b9,
        64'h07b70cf7_16634789,
        64'h873e0347_c783f984,
        64'h3783a451_fef42623,
        64'h47852207_85632781,
        64'hfec42783_fef42623,
        64'h87aa2ac0_00eff984,
        64'h350385be_5f9cf984,
        64'h3783df98_0807071b,
        64'h02faf737_f9843783,
        64'hdc2ff0ef_853e0300,
        64'h05934609_43dcf984,
        64'h3783dfc5_27818b89,
        64'hfe442783_acd9fef4,
        64'h26234785_de6ff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8f984,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_dd4ff0ef,
        64'h853e0300_059343dc,
        64'hf9843783_ae19fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaddaf_e0eff984,
        64'h35036000_0593863e,
        64'h4685fe84_2783fef4,
        64'h242337c5_810007b7,
        64'hc4e19023_47457010,
        64'hd0737010_50730ff0,
        64'h000f818f_f0eff984,
        64'h350385be_863afa04,
        64'h07132781_fe245783,
        64'he7aff0ef_853e4591,
        64'h863afe04_570343dc,
        64'hf9843783_fef41023,
        64'h8ff917fd_6785fe04,
        64'h5703fef4_10230400,
        64'h0793fef4_11234785,
        64'ha65d4785_c2e1ae23,
        64'h4705bf3f_c0ef26e5,
        64'h05130000_15172665,
        64'h85930000_15972040,
        64'h0613a015_14f71363,
        64'h4785873e_0347c783,
        64'hf9843783_c201ae23,
        64'haef94785_c2e1ae23,
        64'h4705c2bf_c0ef2a65,
        64'h05130000_151729e5,
        64'h85930000_15972030,
        64'h0613a015_02f71f63,
        64'h11178793_111117b7,
        64'h873e53dc_f9843783,
        64'hc201ae23_cf91f984,
        64'h3783fc04_3c23fc04,
        64'h3823fc04_3423fc04,
        64'h3023fa04_3c23fa04,
        64'h3823fa04_3423fa04,
        64'h3023f8a4_3c231880,
        64'hf0a2f486_71598082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'hebeff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfc843783_f7eff0ef,
        64'h853e0300_05934609,
        64'h43dcfc84_3783dfc5,
        64'h27818b89_fdc42783,
        64'ha83dfef4_26234785,
        64'hfa2ff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fc84_3783c385,
        64'h27818ff9_67a1fdc4,
        64'h2703fcf4_2e2387aa,
        64'hf90ff0ef_853e0300,
        64'h059343dc_fc843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaf96f,
        64'he0effc84_35036000,
        64'h0593863e_4685fe04,
        64'h27837010_d0737010,
        64'h50730ff0_000ffef4,
        64'h202337c1_010007b7,
        64'hc4e19023_47459d4f,
        64'hf0effc84_350385be,
        64'hfc043603_2781fe64,
        64'h5783835f_f0ef853e,
        64'h4591863a_fe445703,
        64'h43dcfc84_3783fef4,
        64'h12238ff9_17fd6785,
        64'hfe445703_fef41223,
        64'h04000793_fef41323,
        64'h4785fce7_dee303f0,
        64'h07930007_871bfe84,
        64'h2783fef4_24232785,
        64'hfe842783_00078023,
        64'h97bafc04_3703fe84,
        64'h2783aa15_4785c2e1,
        64'hae234705_dd5fc0ef,
        64'h45050513_00001517,
        64'h44858593_00001597,
        64'h1a800613_a835fe04,
        64'h2423c201_ae23a285,
        64'h4785c2e1_ae234705,
        64'he01fc0ef_47c50513,
        64'h00001517_47458593,
        64'h00001597_1a700613,
        64'ha01502f7_19631117,
        64'h87931111_17b7873e,
        64'h53dcfc84_3783c201,
        64'hae23cf91_fc843783,
        64'hfcb43023_fca43423,
        64'h0080f822_fc067139,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aa879f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783939f,
        64'hf0ef853e_03e00593,
        64'h863a9341_1742fe84,
        64'h270343dc_fd843783,
        64'hfef42423_8fd9fe84,
        64'h278357f8_fd843783,
        64'hfef42423_8ff917e1,
        64'h67c1fe84_2703fef4,
        64'h242387aa_93dff0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_04f71963,
        64'h4791873e_57fcfd84,
        64'h3783a15f_f0ef853e,
        64'h02800593_863a0ff7,
        64'h7713fe84_270343dc,
        64'hfd843783_fef42423,
        64'h0027e793_fe842783,
        64'ha039fef4_24230207,
        64'he793fe84_278300f7,
        64'h1963478d_873e0377,
        64'hc783fd84_3783fef4,
        64'h242387aa_a25ff0ef,
        64'h853e0280_059343dc,
        64'hfd843783_93efd0ef,
        64'h3e800513_9f7ff0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe842783,
        64'ha8f5fef4_26234785,
        64'ha1bff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe84,
        64'h2703fef4_242387aa,
        64'ha09ff0ef_853e0300,
        64'h059343dc_fd843783,
        64'haa35fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaa0ff,
        64'he0effd84_35036000,
        64'h0593863e_4681fe44,
        64'h2783fef4_22231007,
        64'h879b03b7_07b7a039,
        64'hfef42223_5007879b,
        64'h03b707b7_00f71963,
        64'h4791873e_57fcfd84,
        64'h3783a02d_fef42223,
        64'h2007879b_03b707b7,
        64'ha825fef4_22236007,
        64'h879b03b7_07b700f7,
        64'h19634791_873e57fc,
        64'hfd843783_02f71763,
        64'h478d873e_0377c783,
        64'hfd843783_02e78ba3,
        64'h4709fd84_3783a031,
        64'h02e78ba3_470dfd84,
        64'h378300f7_186347a1,
        64'h873e4bdc_fd843783,
        64'h00f71f63_4795873e,
        64'h0347c783_fd843783,
        64'h02f71763_4789873e,
        64'h0367c783_fd843783,
        64'ha431fef4_26234785,
        64'h12078c63_2781fec4,
        64'h2783fef4_262387aa,
        64'hae1fe0ef_fd843503,
        64'h60078593_67a1863e,
        64'h4681fe44_2783fef4,
        64'h22230377_c783fd84,
        64'h378302e7_8ba34709,
        64'hfd843783_ac81fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aab23f_e0effd84,
        64'h35037007_8593678d,
        64'h863e4681_4bbcfd84,
        64'h378306f7_1b634785,
        64'h873e0347_c783fd84,
        64'h3783a479_fe042623,
        64'h00e7e563_478d873e,
        64'h4bdcfd84_3783a45d,
        64'h4785c2e1_ae234705,
        64'h900fd0ef_77c50513,
        64'h00001517_77458593,
        64'h00001597_11b00613,
        64'ha01502f7_1e634789,
        64'h873e0367_c783fd84,
        64'h3783c201_ae23acf9,
        64'h4785c2e1_ae234705,
        64'h938fd0ef_7b450513,
        64'h00001517_7ac58593,
        64'h00001597_11a00613,
        64'ha01502f7_1f631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783c201,
        64'hae23cf91_fd843783,
        64'hfca43c23_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aabadf,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfd84,
        64'h3783c6df_f0ef853e,
        64'h03000593_460943dc,
        64'hfd843783_dfc52781,
        64'h8b89fe04_2783a83d,
        64'hfef42623_4785c91f,
        64'hf0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c3852781,
        64'h8ff967a1_fe042703,
        64'hfef42023_87aac7ff,
        64'hf0ef853e_03000593,
        64'h43dcfd84_3783a8bd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_c85fe0ef,
        64'hfd843503_30078593,
        64'h67ad4601_86be2781,
        64'hfe645783_7010d073,
        64'h70105073_0ff0000f,
        64'hc4e19023_4745ebcf,
        64'hf0effd84_350385be,
        64'hfd043603_2781fe64,
        64'h5783d1df_f0ef853e,
        64'h4591863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12238ff9_17fd6785,
        64'hfe445703_fef41223,
        64'h47a1fef4_13234785,
        64'ha201fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aad07f,
        64'he0effd84_35037007,
        64'h8593678d_863e4681,
        64'h4bbcfd84_3783fce7,
        64'hdfe3479d_0007871b,
        64'hfe842783_fef42423,
        64'h2785fe84_27830007,
        64'h802397ba_fd043703,
        64'hfe842783_aaa14785,
        64'hc2e1ae23_4705ae6f,
        64'hd0ef9625_05130000,
        64'h251795a5_85930000,
        64'h25970ba0_0613a835,
        64'hfe042423_c201ae23,
        64'ha2514785_c2e1ae23,
        64'h4705b12f_d0ef98e5,
        64'h05130000_25179865,
        64'h85930000_25970b90,
        64'h0613a015_02f71963,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'hc201ae23_cf91fd84,
        64'h3783fcb4_3823fca4,
        64'h3c231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_e2fff0ef,
        64'h85364591_863e93c1,
        64'h17c28ff9_17fd6785,
        64'hfd645703_43d4fd84,
        64'h3783fef4_26232781,
        64'h87aada9f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783a081,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_e25fe0ef,
        64'hfd843503_6585863e,
        64'h46812781_fd645783,
        64'ha0adfef4_26234785,
        64'ha89d4785_c2e1ae23,
        64'h4705be2f_d0efa5e5,
        64'h05130000_2517a565,
        64'h85930000_259707f0,
        64'h0613a015_c79d2781,
        64'h3037f793_fe842783,
        64'hfef42423_87aae25f,
        64'hf0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_c201ae23,
        64'ha0d94785_c2e1ae23,
        64'h4705c32f_d0efaae5,
        64'h05130000_2517aa65,
        64'h85930000_259707e0,
        64'h0613a015_04f71b63,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'hc201ae23_cf91fd84,
        64'h3783fcf4_1b2387ae,
        64'hfca43c23_1800f022,
        64'hf4067179_80826105,
        64'h644260e2_0001eb7f,
        64'hf0ef853e_85bafea4,
        64'h47039381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef40523,
        64'h87bafef4_05a387b6,
        64'hfef42623_873286ae,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e2853e_87aaea9f,
        64'hf0ef853e_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h05a387ba_fef42623,
        64'h872e87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_0001f63f,
        64'hf0ef853e_85bafe84,
        64'h57039381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef41423,
        64'h87bafef4_05a387b6,
        64'hfef42623_873286ae,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e2853e_87aaf47f,
        64'hf0ef853e_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h05a387ba_fef42623,
        64'h872e87aa_1000e822,
        64'hec061101_80826145,
        64'h74220001_00e79023,
        64'hfd645703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf41b23_87aefca4,
        64'h3c231800_f4227179,
        64'h80826145_74220001,
        64'h00e78023_fd744703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf40ba3,
        64'h87aefca4_3c231800,
        64'hf4227179_80826105,
        64'h6462853e_2781439c,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61056462_853e93c1,
        64'h17c20007_d783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826105,
        64'h6462853e_0ff7f793,
        64'h0007c783_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61616406,
        64'h60a6853e_fec42783,
        64'hfe042623_d3f8fb84,
        64'h37830007_871b0097,
        64'hd79bfd84_2783fcf4,
        64'h2c2302f7_07bbfe04,
        64'h2783fd84_2703fcf4,
        64'h2c2302f7_07bbfdc4,
        64'h27032781_2785fd84,
        64'h2783fcf4_2c238fd9,
        64'hfd842783_0007871b,
        64'h8ff9c007_87936785,
        64'h873e2781_00a7979b,
        64'hfd042783_fcf42c23,
        64'h0167d79b_fcc42783,
        64'hfcf42e23_278100f7,
        64'h17bb4705_27812789,
        64'h27818b9d_27810077,
        64'hd79bfcc4_2783fef4,
        64'h20232781_00f717bb,
        64'h47052781_8bbd2781,
        64'h0087d79b_fd042783,
        64'h02e78aa3_fb843783,
        64'h0ff7f713_8bbd0ff7,
        64'hf7932781_0127d79b,
        64'hfd442783_fcf42a23,
        64'h278187aa_a11fd0ef,
        64'h853e9381_17822781,
        64'h27f143dc_fb843783,
        64'hfcf42823_278187aa,
        64'ha2dfd0ef_853e9381,
        64'h17822781_27e143dc,
        64'hfb843783_fcf42623,
        64'h278187aa_a49fd0ef,
        64'h853e9381_17822781,
        64'h27d143dc_fb843783,
        64'hfcf42423_278187aa,
        64'ha65fd0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_a23dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa9e2f_f0effb84,
        64'h35039007_85936785,
        64'h863e4681_4bbcfb84,
        64'h3783aab1_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'ha10ff0ef_fb843503,
        64'h30000593_863e4681,
        64'h4bbcfb84_3783cbb8,
        64'h12340737_fb843783,
        64'hc7f8fb84_37830007,
        64'h871b87aa_b85fd0ef,
        64'h853e45f1_43dcfb84,
        64'h3783c7b8_fb843783,
        64'h0007871b_87aab9ff,
        64'hd0ef853e_45e143dc,
        64'hfb843783_c3f8fb84,
        64'h37830007_871b87aa,
        64'hbb9fd0ef_853e45d1,
        64'h43dcfb84_3783c3b8,
        64'hfb843783_0007871b,
        64'h87aabd3f_d0ef853e,
        64'h45c143dc_fb843783,
        64'haaedfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaaaef,
        64'hf0effb84_35032000,
        64'h05934601_4681db98,
        64'h4705fb84_3783c789,
        64'h27818ff9_400007b7,
        64'hfe842703_fa07dde3,
        64'hfe842783_fef42423,
        64'h87aab8ff_d0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783aca1,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_b0cff0ef,
        64'hfb843503_10000593,
        64'h40ff8637_4681a091,
        64'hfe042423_a459fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aab3af_f0effb84,
        64'h35034581_46014681,
        64'ha46dfef4_26234785,
        64'he7892781_8ff967c1,
        64'hfe442703_fef42223,
        64'h87aac0ff_d0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fb843783,
        64'hcb8d47dc_fb843783,
        64'h02f70e63_400007b7,
        64'h873e2781_8ff9c000,
        64'h07b7873e_579cfb84,
        64'h3783a601_4785c2e1,
        64'hae234705_93dfd0ef,
        64'hf9850513_00002517,
        64'hf9858593_00002597,
        64'h68900613_a01504f7,
        64'h11634789_873e0367,
        64'hc783fb84_3783c201,
        64'hae23ae25_4785c2e1,
        64'hae234705_975fd0ef,
        64'hfd050513_00002517,
        64'hfd058593_00002597,
        64'h68800613_a01502f7,
        64'h1f631117_87931111,
        64'h17b7873e_53dcfb84,
        64'h3783c201_ae23cf91,
        64'hfb843783_faa43c23,
        64'h0880e0a2_e486715d,
        64'h80826121_744270e2,
        64'h00017010_d0737010,
        64'h50730ff0_000fd55f,
        64'hd0ef853a_85be2781,
        64'h08078793_fd843783,
        64'h93010207_97132781,
        64'h0587879b_43dcfd84,
        64'h378300e7_912397b6,
        64'h078e07c1_93810206,
        64'h1793fd84_36839341,
        64'h03079713_02f707bb,
        64'h0006861b_36fdfec4,
        64'h268393c1_17c2fe44,
        64'h27839341_03079713,
        64'hfd442783_00e79023,
        64'h02300713_97ba078e,
        64'h07c19381_1782fd84,
        64'h37032781_37fdfec4,
        64'h2783c3d8_97b6078e,
        64'h07c19381_02061793,
        64'hfd843683_0007871b,
        64'h9fb90006_861b36fd,
        64'hfec42683_27810107,
        64'h979bfe84_27830007,
        64'h871bfc84_3783f8e7,
        64'hebe32781_fe842783,
        64'h0007871b_37fdfec4,
        64'h2783fef4_24232785,
        64'hfe842783_00079123,
        64'h97ba078e_07c1fe84,
        64'h6783fd84_370300e7,
        64'h90230210_071397ba,
        64'h078e07c1_fe846783,
        64'hfd843703_c3d897b6,
        64'h078e07c1_fe846783,
        64'hfd843683_0007871b,
        64'h9fb92781_0107979b,
        64'hfe842783_0007871b,
        64'hfc843783_a8b1fe04,
        64'h2423fef4_26232785,
        64'hfec42783_c7912781,
        64'h8ff917fd_67c1873e,
        64'h278102f7_07bbfe44,
        64'h2783fd44_2703fef4,
        64'h26230107_d79b2781,
        64'h02f707bb_fe442783,
        64'hfd442703_a835fef4,
        64'h26234785_00f77663,
        64'h67c1873e_278102f7,
        64'h07bbfe44_2783fd44,
        64'h2703fef4_22238ff9,
        64'h17fd6785_fe442703,
        64'hfef42223_87aaf0ff,
        64'hd0ef853e_459143dc,
        64'hfd843783_fe042223,
        64'hfe042423_fe042623,
        64'hfcf42a23_fcc43423,
        64'h87aefca4_3c230080,
        64'hf822fc06_71398082,
        64'h61457402_70a2853e,
        64'hfec42783_0001a011,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_e1cff0ef,
        64'hfd843503_70000593,
        64'h863e4681_4bbcfd84,
        64'h3783fe04_2623fca4,
        64'h3c231800_f022f406,
        64'h71798082_61217442,
        64'h70e2853e_fec42783,
        64'hfe042623_fd7fd0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe442783,
        64'ha00dfef4_26234785,
        64'hffbfd0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe44,
        64'h2703fef4_222387aa,
        64'hfe9fd0ef_853e0300,
        64'h059343dc_fd843783,
        64'ha08dfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaec6f,
        64'hf0effd84_35039007,
        64'h85936789_863e86ba,
        64'hfd442783_fd042703,
        64'hc4e19023_02700713,
        64'ha869fef4_26234785,
        64'hc3a92781_fec42783,
        64'hfef42623_87aaefef,
        64'hf0effd84_35038007,
        64'h85936789_863e86ba,
        64'hfd442783_fd042703,
        64'hc4e19023_470d02f7,
        64'h1d634785_0007871b,
        64'hfd042783_7010d073,
        64'h70105073_0ff0000f,
        64'h146000ef_fd843503,
        64'h85befc84_3603fd04,
        64'h2783a8f5_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h081000ef_fd843503,
        64'h20000593_02f70363,
        64'h20000793_873e2781,
        64'h87aa826f_e0ef853e,
        64'h93811782_27812791,
        64'h43dcfd84_3783a281,
        64'hfef42623_4785e789,
        64'h27818ff9_67c1fe84,
        64'h2703fef4_242387aa,
        64'h854fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783cb8d,
        64'h47dcfd84_378302f7,
        64'h0e634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_fd843783,
        64'h00f71f63_4789873e,
        64'h0367c783_fd843783,
        64'hfcf42823_87bafcf4,
        64'h2a23fcd4_34238732,
        64'h87aefca4_3c230080,
        64'hf822fc06_71398082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'h8d4fe0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_9befe0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe442783,
        64'ha83dfef4_26234785,
        64'h9e2fe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe44,
        64'h2703fef4_222387aa,
        64'h9d0fe0ef_853e0300,
        64'h059343dc_fd843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa8aff,
        64'hf0effd84_35032007,
        64'h85936785_863e86ba,
        64'hfd442783_fd042703,
        64'hc4e19023_03700713,
        64'ha85dfef4_26234785,
        64'hc3a92781_fec42783,
        64'hfef42623_87aa8e7f,
        64'hf0effd84_35031007,
        64'h85936785_863e86ba,
        64'hfd442783_fd042703,
        64'hc4e19023_474d02f7,
        64'h1d634785_0007871b,
        64'hfd042783_7010d073,
        64'h70105073_0ff0000f,
        64'h32e000ef_fd843503,
        64'h85befc84_3603fd04,
        64'h2783aa21_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h269000ef_fd843503,
        64'h20000593_02f70363,
        64'h20000793_873e2781,
        64'h87aaa0ef_e0ef853e,
        64'h93811782_27812791,
        64'h43dcfd84_3783aab1,
        64'hfef42623_4785e789,
        64'h27818ff9_67c1fe84,
        64'h2703fef4_242387aa,
        64'ha3cfe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783cb8d,
        64'h47dcfd84_378302f7,
        64'h0e634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_fd843783,
        64'h00f71f63_4789873e,
        64'h0367c783_fd843783,
        64'hfcf42823_87bafcf4,
        64'h2a23fcd4_34238732,
        64'h87aefca4_3c230080,
        64'hf822fc06_71398082,
        64'h61457422_853efec4,
        64'h27830001_a0110001,
        64'ha0210001_a031fef4,
        64'h26238fd9_fd442783,
        64'hfec42703_a831fef4,
        64'h262301a7_e793fec4,
        64'h2783a02d_fef42623,
        64'h03a7e793_fec42783,
        64'ha825fef4_262301a7,
        64'he793fec4_2783a099,
        64'hfef42623_0027e793,
        64'hfec42783_a891fef4,
        64'h262303a7_e793fec4,
        64'h2783a08d_fef42623,
        64'h03a7e793_fec42783,
        64'ha885fef4_262301a7,
        64'he793fec4_2783a8bd,
        64'hfef42623_0097e793,
        64'hfec42783_a071fef4,
        64'h262303a7_e793fec4,
        64'h2783a869_fef42623,
        64'h01a7e793_fec42783,
        64'h00f71963_4785873e,
        64'h0347c783_fd843783,
        64'ha865fef4_262301a7,
        64'he793fec4_2783a0d9,
        64'hfef42623_01a7e793,
        64'hfec42783_a8d1fef4,
        64'h262301b7_e793fec4,
        64'h2783a0cd_fef42623,
        64'h03a7e793_fec42783,
        64'h00f71963_4785873e,
        64'h0347c783_fd843783,
        64'ha201fef4_262301b7,
        64'he793fec4_2783a239,
        64'hfef42623_01b7e793,
        64'hfec42783_aa31fef4,
        64'h26230097_e793fec4,
        64'h2783a22d_fef42623,
        64'h0027e793_fec42783,
        64'haa390ef7_05639007,
        64'h879367ad_0007871b,
        64'h10e68a63_30070713,
        64'h672d0007_869b10e6,
        64'h8a63a007_0713672d,
        64'h0007869b_a2a916f7,
        64'h0363a007_87936791,
        64'h0007871b_0ee68d63,
        64'hd0070713_67250007,
        64'h869b0ae6_89636007,
        64'h07136721_0007869b,
        64'h02d76863_70070713,
        64'h67250007_869b14e6,
        64'h80637007_07136725,
        64'h0007869b_aa4914f7,
        64'h08638007_87936789,
        64'h0007871b_18e68b63,
        64'h40070713_670d0007,
        64'h869b16e6_86639007,
        64'h07136709_0007869b,
        64'haa7d16f7_07632007,
        64'h87936785_0007871b,
        64'h16e68e63_50070713,
        64'h67050007_869b18e6,
        64'h85633007_07136705,
        64'h0007869b_02d76863,
        64'h70070713_67050007,
        64'h869b1ae6_8a637007,
        64'h07136705_0007869b,
        64'h06d76c63_70070713,
        64'h670d0007_869b20e6,
        64'h84637007_0713670d,
        64'h0007869b_a40d1cf7,
        64'h0263b007_87936785,
        64'h0007871b_1ce68963,
        64'h67050007_869b1ce6,
        64'h8e63c007_07136705,
        64'h0007869b_a4a91af7,
        64'h02637000_07930007,
        64'h871b1ee6_85639007,
        64'h07136705_0007869b,
        64'h1c070663_27018007,
        64'h871b02d7_6563a007,
        64'h07136705_0007869b,
        64'h20e68f63_a0070713,
        64'h67050007_869ba471,
        64'h18f70863_30000793,
        64'h0007871b_1ae68563,
        64'h50000713_0007869b,
        64'h2ae68e63_40000713,
        64'h0007869b_ac4d18f7,
        64'h0d631000_07930007,
        64'h871b2c07_09630007,
        64'h871b00d7_6d632000,
        64'h07130007_869b1ce6,
        64'h84632000_07130007,
        64'h869b04d7_6c636000,
        64'h07130007_869b20e6,
        64'h85636000_07130007,
        64'h869b0cd7_6d631007,
        64'h07136705_0007869b,
        64'h2ae68a63_10070713,
        64'h67050007_869bfd44,
        64'h2783fef4_2623fd44,
        64'h2783fcf4_2a2387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61217442,
        64'h70e2853e_fec42783,
        64'hfe042623_edefe0ef,
        64'h853e0300_05934605,
        64'h43dcfd84_3783d3a9,
        64'h27818b85_fe042783,
        64'ha00defcf_e0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hfef42623_4789e781,
        64'h27819bf9_fec42783,
        64'hfef42623_87aaeeef,
        64'he0ef853e_03200593,
        64'h43dcfd84_3783c3a1,
        64'h27818ff9_67a1fe04,
        64'h2703a899_f46fe0ef,
        64'h853e0300_05930200,
        64'h061343dc_fd843783,
        64'hcf812781_0207f793,
        64'h278187aa_f2cfe0ef,
        64'h853e0300_059343dc,
        64'hfd843783_02f71b63,
        64'h30078793_67850007,
        64'h871bfd44_278300f7,
        64'h0b635007_87936785,
        64'h0007871b_fd442783,
        64'hfef42023_87aaf66f,
        64'he0ef853e_03000593,
        64'h43dcfd84_3783f4cf,
        64'he0ef853a_85be2781,
        64'h8fd52781_c401d783,
        64'h0007869b_0107979b,
        64'hfe442783_93010207,
        64'h97132781_27b143dc,
        64'hfd843783_a219fef4,
        64'h26234785_c7892781,
        64'h0207f793_fe442783,
        64'hcb992781_8b89fe84,
        64'h2783fef4_242387aa,
        64'hf2cfe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_378302f7,
        64'h0f633007_87936785,
        64'h0007871b_fd442783,
        64'h04f70863_50078793,
        64'h67850007_871bfd44,
        64'h2783fef4_22238ff9,
        64'h17fd6791_fe442703,
        64'hfef42223_87aa1880,
        64'h00effd84_350385be,
        64'hfd442783_85ffe0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783875f_e0ef853a,
        64'h03000593_fff78613,
        64'h67c143d8_fd843783,
        64'h827fe0ef_853e85ba,
        64'hfd042703_93811782,
        64'h278127a1_43dcfd84,
        64'h3783925f_e0ef853e,
        64'h02e00593_463943dc,
        64'hfd843783_8b7fe0ef,
        64'h853e4599_863a9341,
        64'h1742fcc4_270343dc,
        64'hfd843783_aaddfef4,
        64'h26234785_a4094785,
        64'hc2e1ae23_4705cf6f,
        64'he0efb525_05130000,
        64'h3517b525_85930000,
        64'h359744c0_0613a015,
        64'hc79d2781_8b85fe84,
        64'h2783fef4_242387aa,
        64'h835fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783c201,
        64'hae23ac81_4785c2e1,
        64'hae234705_d44fe0ef,
        64'hba050513_00003517,
        64'hba058593_00003597,
        64'h44b00613_a01504f7,
        64'h1a631117_87931111,
        64'h17b7873e_53dcfd84,
        64'h3783c201_ae23cf91,
        64'hfd843783_fcf42623,
        64'h87bafcf4_282387b2,
        64'hfcf42a23_873687ae,
        64'hfca43c23_0080f822,
        64'hfc067139_80826145,
        64'h740270a2_853efec4,
        64'h27830001_fcf719e3,
        64'h01f007b7_873e2781,
        64'h8ff901f0_07b7fe84,
        64'h2703fef4_242387aa,
        64'h8ddfe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783a839,
        64'hfef42423_87aa8fbf,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_80ffe0ef,
        64'h3e800513_9effe0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0047e793,
        64'h93c117c2_fe442783,
        64'h43d8fd84_3783fef4,
        64'h222387aa_9ddfe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_d3ed2781,
        64'h8b89fe44_2783fef4,
        64'h222387aa_9fdfe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a821fef4,
        64'h222387aa_a15fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a5ffe0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0017e793,
        64'h93c117c2_fe442783,
        64'h43d8fd84_3783fef4,
        64'h222387aa_a4dfe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a211fef4,
        64'h26234785_e7892781,
        64'h8ba12781_fe245783,
        64'hfef41123_87aaa77f,
        64'he0ef853e_03e00593,
        64'h43dcfd84_37838e9f,
        64'he0ef3887_85136785,
        64'hacbfe0ef_853e03e0,
        64'h0593863a_fe245703,
        64'h43dcfd84_3783fef4,
        64'h11230087_e793fe24,
        64'h5783fef4_112387aa,
        64'hab9fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'hb03fe0ef_853e02c0,
        64'h0593863a_fe245703,
        64'h43dcfd84_3783fef4,
        64'h11239be9_fe245783,
        64'hfef41123_87aaaeff,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783ffe1,
        64'h27818ff9_01f007b7,
        64'hfe842703_fef42423,
        64'h87aaa77f_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'ha839fef4_242387aa,
        64'ha95fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783fef4,
        64'h26234785_c7812781,
        64'hfec42783_fef42623,
        64'h87aa2120_00effd84,
        64'h3503b007_85936785,
        64'h46014681_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623f3e5_27818b89,
        64'h2781feb4_4783fef4,
        64'h05a387aa_c1dfe0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_a821fef4,
        64'h05a387aa_c35fe0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_c7ffe0ef,
        64'h853e02f0_05934609,
        64'h43dcfd84_3783c11f,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c27fe0ef,
        64'h853a0300_0593fff7,
        64'h861367c1_43d8fd84,
        64'h378302e7_8a234709,
        64'hfd843783_a03102e7,
        64'h8a234705_fd843783,
        64'hc7992781_fec42783,
        64'hfef42623_87aa2de0,
        64'h00effd84_35031000,
        64'h059340ff_86374681,
        64'ha855fef4_26234785,
        64'ha0c14785_c2e1ae23,
        64'h470589bf_e0efef65,
        64'h05130000_3517ef65,
        64'h85930000_35973ac0,
        64'h0613a015_c79d2781,
        64'hfec42783_fef42623,
        64'h87aa32a0_00effd84,
        64'h35034581_46014681,
        64'hae3fe0ef_71078513,
        64'h6789c201_ae23a239,
        64'h4785c2e1_ae234705,
        64'h8e9fe0ef_f4450513,
        64'h00003517_f4458593,
        64'h00003597_3ab00613,
        64'ha01504f7_1a631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783c201,
        64'hae23cf91_fd843783,
        64'hfca43c23_1800f022,
        64'hf4067179_8082614d,
        64'h64ea740a_70aa853e,
        64'hfdc42783_0001a011,
        64'h0001a021_0001a031,
        64'hfcf42e23_4785cb89,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_4e4010ef,
        64'hf5843503_20000593,
        64'h02f71763_4785873e,
        64'h0347c783_f5843783,
        64'h00f71a63_4791873e,
        64'h57fcf584_37830001,
        64'ha0b9fcf4_2e234785,
        64'hc7912781_fdc42783,
        64'hfcf42e23_87aa71e0,
        64'h20eff584_350385be,
        64'hfd442783_fcf42a23,
        64'h1007879b_03a207b7,
        64'heb950a27_c7830ae7,
        64'h87931ffe_d797a071,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_065010ef,
        64'hf5843503_02f71163,
        64'h4791873e_57fcf584,
        64'h3783a865_fcf42e23,
        64'h478500f7_06634785,
        64'h873e0b97_c7830f67,
        64'h87931ffe_d79704f7,
        64'h16634791_873e57fc,
        64'hf5843783_00f70963,
        64'h4795873e_57fcf584,
        64'h3783a8c5_fcf42e23,
        64'h478500f7_06634789,
        64'h873e0b97_c78312e7,
        64'h87931ffe_d79702f7,
        64'h1063479d_873e57fc,
        64'hf5843783_aa29fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa6340_20eff584,
        64'h35031625_85931ffe,
        64'hd597a281_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h607010ef_f5843503,
        64'h0cf70b63_4799873e,
        64'h57fcf584_3783d7f8,
        64'h4719f584_3783a029,
        64'hd7f84715_f5843783,
        64'h00e7f763_4785873e,
        64'h0377c783_f5843783,
        64'hcf912781_8b892781,
        64'h0c47c783_1c478793,
        64'h1ffed797_a825d7f8,
        64'h4711f584_378300e7,
        64'hf7634785_873e0377,
        64'hc783f584_3783cf91,
        64'h27818bb1_27810c47,
        64'hc7831f27_87931ffe,
        64'hd797a09d_d7f8471d,
        64'hf5843783_00e7f763,
        64'h4785873e_0377c783,
        64'hf5843783_cf912781,
        64'h0307f793_27810c47,
        64'hc7832227_87931ffe,
        64'hd797d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0d47c783_23c78793,
        64'h1ffed797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0087979b_27810d57,
        64'hc7832627_87931ffe,
        64'hd79753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810107,
        64'h979b2781_0d67c783,
        64'h28878793_1ffed797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h0187979b_27810d77,
        64'hc7832aa7_87931ffe,
        64'hd797a461_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h7a2020ef_f5843503,
        64'h2d058593_1ffed597,
        64'ha47dfcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa2870,
        64'h10eff584_350328f7,
        64'h12634795_873e0347,
        64'hc783f584_3783acf1,
        64'hfcf42e23_478528f7,
        64'h0d634785_873e0b97,
        64'hc78331a7_87931ffe,
        64'hd797ace5_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h013020ef_f5843503,
        64'h34058593_1ffed597,
        64'hae39fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa7e50,
        64'h10eff584_3503d7f8,
        64'h4715f584_37832ee7,
        64'hfd634785_873e0377,
        64'hc783f584_37833007,
        64'h85632781_8b892781,
        64'h0c47c783_38c78793,
        64'h1ffed797_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810d47_c7833a67,
        64'h87931ffe_d79753f8,
        64'hf5843783_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810087_979b2781,
        64'h0d57c783_3cc78793,
        64'h1ffed797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0107979b_27810d67,
        64'hc7833f27_87931ffe,
        64'hd79753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b0187_979b2781,
        64'h0d77c783_41478793,
        64'h1ffed797_aecdfcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa10d0_20eff584,
        64'h350343a5_85931ffe,
        64'hd597a921_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h3f1010ef_f5843503,
        64'h14f71f63_4785873e,
        64'h0367c783_f5843783,
        64'h16e7f763_478d873e,
        64'h0357c783_f5843783,
        64'h16f71f63_4789873e,
        64'h0347c783_f5843783,
        64'ha19dfcf4_2e234785,
        64'h42078363_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h12e020ef_f5843503,
        64'hd7f84715_f5843783,
        64'h44e7f363_4785873e,
        64'h0377c783_f5843783,
        64'h44078b63_27818b89,
        64'h2781f9d4_47834607,
        64'h82630004_c78302e7,
        64'h8e234705_f5843783,
        64'h80aff0ef_3e800513,
        64'h9eaff0ef_853a02c0,
        64'h0593863e_93c117c2,
        64'h0047e793_fda45783,
        64'h43d8f584_3783fcf4,
        64'h1d2387aa_9d4ff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_d3e52781,
        64'h8b892781_fda45783,
        64'hfcf41d23_87aa9f6f,
        64'hf0ef853e_02c00593,
        64'h43dcf584_3783a821,
        64'hfcf41d23_87aaa0ef,
        64'hf0ef853e_02c00593,
        64'h43dcf584_3783a58f,
        64'hf0ef853a_02c00593,
        64'h863e93c1_17c20017,
        64'he793fda4_578343d8,
        64'hf5843783_fcf41d23,
        64'h87aaa42f_f0ef853e,
        64'h02c00593_43dcf584,
        64'h3783a3a5_fcf42e23,
        64'h4785e789_27818ba1,
        64'h2781fd24_5783fcf4,
        64'h192387aa_a6cff0ef,
        64'h853e03e0_059343dc,
        64'hf5843783_8deff0ef,
        64'h38878513_6785ac0f,
        64'hf0ef853e_03e00593,
        64'h863afd24_570343dc,
        64'hf5843783_fcf41923,
        64'h0087e793_fd245783,
        64'hfcf41923_87aaaaef,
        64'hf0ef853e_03e00593,
        64'h43dcf584_3783af8f,
        64'hf0ef853e_02c00593,
        64'h863afd24_570343dc,
        64'hf5843783_fcf41923,
        64'h9be9fd24_5783fcf4,
        64'h192387aa_ae4ff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_14079d63,
        64'h03c7c783_f5843783,
        64'h16f71363_47a1873e,
        64'h4bdcf584_378316e7,
        64'hfa63478d_873ef9d4,
        64'h47831807_d0634187,
        64'hd79b0187_979b0024,
        64'hc7836207_9e632781,
        64'hfdc42783_fcf42e23,
        64'h87aa1460_20eff584,
        64'h350385be_f9040793,
        64'hadb9fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa6370,
        64'h10eff584_3503c385,
        64'h27818b91_27810014,
        64'hc783a561_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h483010ef_f5843503,
        64'h85a6a565_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h2e5020ef_f5843503,
        64'h26f71263_4785873e,
        64'h0347c783_f5843783,
        64'hadd9fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa4500,
        64'h10eff584_3503add5,
        64'hfcf42e23_4785adf5,
        64'hfcf42e23_4785cb89,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_017020ef,
        64'hf5843503_85be5f9c,
        64'hf5843783_df98a807,
        64'h071b018c_c737f584,
        64'h3783af05_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h6cc010ef_f5843503,
        64'h04f71b63_4795873e,
        64'h0347c783_f5843783,
        64'h00f70a63_4789873e,
        64'h0347c783_f5843783,
        64'ha7bdfcf4_2e234785,
        64'hc3d12781_fdc42783,
        64'hfcf42e23_87aa0890,
        64'h20eff584_350385be,
        64'h5f9cf584_3783df98,
        64'h8407071b_017d8737,
        64'hf5843783_a801df98,
        64'hac07071b_0121f737,
        64'hf5843783_00f71a63,
        64'h4789873e_0367c783,
        64'hf5843783_7c40006f,
        64'hfcf42e23_4785c791,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_935ff0ef,
        64'hf5843503_06f71c63,
        64'h4785873e_0347c783,
        64'hf5843783_7f40006f,
        64'hfcf42e23_478500f7,
        64'h07634795_873e0347,
        64'hc783f584_378300f7,
        64'h0f634789_873e0347,
        64'hc783f584_378302f7,
        64'h07634785_873e0347,
        64'hc783f584_378302f7,
        64'h02e34785_0007871b,
        64'hfdc42783_fcf42e23,
        64'h87aa0530_00eff584,
        64'h3503a839_02e78a23,
        64'h4715f584_378300f7,
        64'h18634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_f5843783,
        64'h0750006f_4785c2e1,
        64'hae234705_9b4ff0ef,
        64'h81050513_00004517,
        64'h81058593_00004597,
        64'h24000613_a01d04f7,
        64'h18634789_873e0367,
        64'hc783f584_3783df98,
        64'ha807071b_00062737,
        64'hf5843783_02078e23,
        64'hf5843783_02e78a23,
        64'h4705f584_378302e7,
        64'h8ba34705_f5843783,
        64'hc201ae23_0d90006f,
        64'h4785c2e1_ae234705,
        64'ha18ff0ef_87450513,
        64'h00004517_87458593,
        64'h00004597_23f00613,
        64'ha01d06f7_15631117,
        64'h87931111_17b7873e,
        64'h53dcf584_3783c201,
        64'hae23cf91_f5843783,
        64'hfc043423_fc043023,
        64'hfa043c23_fa043823,
        64'hfa043423_fa043023,
        64'hf8043c23_f8043823,
        64'h0004b023_00579493,
        64'h839507fd_f8078793,
        64'hfe040793_f4a43c23,
        64'h1900ed26_f122f506,
        64'h71718082_61616406,
        64'h60a6853e_fec42783,
        64'hfe042623_d3f8fb84,
        64'h37830007_871b00a7,
        64'h979b2781_27852781,
        64'h8ff917fd_004007b7,
        64'h873e2781_0087d79b,
        64'hfc442783_02f71663,
        64'h4785873e_27818b8d,
        64'h27810167_d79bfcc4,
        64'h2783a081_d3f8fb84,
        64'h37830007_871b0097,
        64'hd79bfd04_2783fcf4,
        64'h282302f7_07bbfd84,
        64'h2783fd04_2703fcf4,
        64'h282302f7_07bbfd44,
        64'h27032781_2785fd04,
        64'h2783fcf4_28238fd9,
        64'hfd042783_0007871b,
        64'h8ff9c007_87936785,
        64'h873e2781_00a7979b,
        64'hfc842783_fcf42823,
        64'h0167d79b_fc442783,
        64'hfcf42a23_278100f7,
        64'h17bb4705_27812789,
        64'h27818b9d_27810077,
        64'hd79bfc44_2783fcf4,
        64'h2c232781_00f717bb,
        64'h47052781_8bbd2781,
        64'h0087d79b_fc842783,
        64'he3c52781_8b8d2781,
        64'h0167d79b_fcc42783,
        64'hfcf42623_278187aa,
        64'heacff0ef_853e9381,
        64'h17822781_27f143dc,
        64'hfb843783_fcf42423,
        64'h278187aa_ec8ff0ef,
        64'h853e9381_17822781,
        64'h27e143dc_fb843783,
        64'hfcf42223_278187aa,
        64'hee4ff0ef_853e9381,
        64'h17822781_27d143dc,
        64'hfb843783_fcf42023,
        64'h278187aa_f00ff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'ha28dfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa67f0,
        64'h00effb84_35039007,
        64'h85936785_863e4681,
        64'h4bbcfb84_3783d7d5,
        64'h4bbcfb84_3783cbb8,
        64'hfb843783_0007871b,
        64'h8ff977c1_873e2781,
        64'h87aaf5ef_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783a2c1,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_6dd000ef,
        64'hfb843503_30000593,
        64'h46014681_c7f8fb84,
        64'h37830007_871b87aa,
        64'h841ff0ef_853e45f1,
        64'h43dcfb84_3783c7b8,
        64'hfb843783_0007871b,
        64'h87aa85bf_f0ef853e,
        64'h45e143dc_fb843783,
        64'hc3f8fb84_37830007,
        64'h871b87aa_875ff0ef,
        64'h853e45d1_43dcfb84,
        64'h3783c3b8_fb843783,
        64'h0007871b_87aa88ff,
        64'hf0ef853e_45c143dc,
        64'hfb843783_a4b9fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa76b0_00effb84,
        64'h35032000_05934601,
        64'h4681ac95_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h565000ef_fb843503,
        64'h02e78e23_4705fb84,
        64'h3783c78d_27818ff9,
        64'h010007b7_fe842703,
        64'hdb984705_fb843783,
        64'hc7892781_8ff94000,
        64'h07b7fe84_2703f407,
        64'hdde3fe84_2783fef4,
        64'h242387aa_881ff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'ha4cdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa7ff0,
        64'h00effb84_35039007,
        64'h859367ad_863e4681,
        64'hfe442783_fef42223,
        64'h8fd90100_07b7fe44,
        64'h270300f7_196347a1,
        64'h873e4bdc_fb843783,
        64'h02f71063_4789873e,
        64'h0367c783_fb843783,
        64'hfef42223_40ff87b7,
        64'ha689fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa05e0,
        64'h10effb84_35037007,
        64'h8593678d_46014681,
        64'ha055fe04_242302e7,
        64'h8aa34709_fb843783,
        64'ha03102e7_8aa34705,
        64'hfb843783_00f70863,
        64'h1aa00793_0007871b,
        64'hfe842783_fef42423,
        64'h87aa94ff_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783f3e5,
        64'h27818b89_2781fe34,
        64'h4783fef4_01a387aa,
        64'ha91ff0ef_853e02f0,
        64'h059343dc_fb843783,
        64'ha821fef4_01a387aa,
        64'haa9ff0ef_853e02f0,
        64'h059343dc_fb843783,
        64'haf3ff0ef_853e02f0,
        64'h05934609_43dcfb84,
        64'h378304f7_18634789,
        64'h0007871b_fec42783,
        64'ha129fef4_26234785,
        64'h00f70663_47890007,
        64'h871bfec4_2783cf81,
        64'h2781fec4_2783fef4,
        64'h262387aa_134010ef,
        64'hfb843503_80078593,
        64'h67851aa0_06134681,
        64'ha189fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa15e0,
        64'h10effb84_35034581,
        64'h46014681_a19dfef4,
        64'h26234785_e7892781,
        64'h8ff967c1_fdc42703,
        64'hfcf42e23_87aaa33f,
        64'hf0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfb843783_cb8d47dc,
        64'hfb843783_02f70e63,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cfb84_3783a975,
        64'h4785c2e1_ae234705,
        64'hf60ff0ef_dbc50513,
        64'h00004517_dbc58593,
        64'h00004597_16200613,
        64'ha01504f7_11634789,
        64'h873e0367_c783fb84,
        64'h3783cbd8_4711fb84,
        64'h3783c201_ae23a9f5,
        64'h4785c2e1_ae234705,
        64'hfa0ff0ef_dfc50513,
        64'h00004517_dfc58593,
        64'h00004597_16100613,
        64'ha01504f7_13631117,
        64'h87931111_17b7873e,
        64'h53dcfb84_3783c201,
        64'hae23cf91_fb843783,
        64'hfaa43c23_0880e0a2,
        64'he486715d_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623be1f,
        64'hf0ef853e_45912000,
        64'h061343dc_fd843783,
        64'hc4e19023_474dbf9f,
        64'hf0ef853e_03a00593,
        64'h460143dc_fd843783,
        64'hc0bff0ef_853e0380,
        64'h05934601_43dcfd84,
        64'h3783c1df_f0ef853a,
        64'h03600593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hc33ff0ef_853a0340,
        64'h0593eff7_861367c1,
        64'h43d8fd84_3783cc9f,
        64'hf0ef853e_02800593,
        64'h464143dc_fd843783,
        64'hcdbff0ef_853a0290,
        64'h0593863e_0ff7f793,
        64'h0017e793_feb44783,
        64'h43d8fd84_3783fe04,
        64'h05a3a019_fef405a3,
        64'h47a9c789_27818ff9,
        64'h040007b7_873e579c,
        64'hfd843783_a005fef4,
        64'h05a347b1_c7892781,
        64'h8ff90200_07b7873e,
        64'h579cfd84_3783a82d,
        64'hfef405a3_47b9c789,
        64'h27818ff9_010007b7,
        64'h873e579c_fd843783,
        64'ha8c5fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa0c00,
        64'h30effd84_3503a807,
        64'h85930006_27b7b19f,
        64'hf0ef0c80_051300f7,
        64'h16634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_fd843783,
        64'h02f71363_4789873e,
        64'h0367c783_fd843783,
        64'hda3ff0ef_853e0290,
        64'h0593463d_43dcfd84,
        64'h3783a811_db7ff0ef,
        64'h853e0290_0593463d,
        64'h43dcfd84_378300f7,
        64'h1c634789_873e0367,
        64'hc783fd84_3783d798,
        64'hfd843783_0007871b,
        64'h87aac8ff_f0ef853e,
        64'h93811782_27810407,
        64'h879b43dc_fd843783,
        64'h02e78b23_fd843783,
        64'h0ff7f713_87aad4ff,
        64'hf0ef853e_0fe00593,
        64'h43dcfd84_3783f3e5,
        64'h27818b85_2781fea4,
        64'h4783fef4_052387aa,
        64'hdf1ff0ef_853e02f0,
        64'h059343dc_fd843783,
        64'ha821fef4_052387aa,
        64'he09ff0ef_853e02f0,
        64'h059343dc_fd843783,
        64'he53ff0ef_853e02f0,
        64'h05934605_43dcfd84,
        64'h3783c0df_f0ef3e80,
        64'h0513e6df_f0ef853e,
        64'h02900593_460143dc,
        64'hfd843783_a811e81f,
        64'hf0ef853e_02900593,
        64'h464143dc_fd843783,
        64'hac354785_c2e1ae23,
        64'h4705a33f_f0ef08e5,
        64'h05130000_451708e5,
        64'h85930000_45970b50,
        64'h0613a015_02f71e63,
        64'h4789873e_27810ff7,
        64'hf7932781_87aae0ff,
        64'hf0ef853e_0fe00593,
        64'h43dcfd84_37830607,
        64'hb823fd84_3783d7f8,
        64'h4719fd84_37830607,
        64'ha223fd84_378302e7,
        64'h8023fd84_37830207,
        64'hc703fd04_3783cfd8,
        64'hfd843783_4fd8fd04,
        64'h3783cf98_fd843783,
        64'h4f98fd04_3783cbd8,
        64'hfd843783_4bd8fd04,
        64'h3783cb98_fd843783,
        64'h4b98fd04_3783c7d8,
        64'hfd843783_47d8fd04,
        64'h3783d3d8_1117071b,
        64'h11111737_fd843783,
        64'hc798fd84_37834798,
        64'hfd043783_c3d8fcc4,
        64'h2703fd84_378300e7,
        64'h9023fd84_37830007,
        64'hd703fd04_3783c201,
        64'hae23ae39_4785c2e1,
        64'hae234705_b15ff0ef,
        64'h17050513_00004517,
        64'h17058593_00004597,
        64'h0b400613_a015c3fd,
        64'hfd043783_c201ae23,
        64'hc799fd84_3783fcf4,
        64'h262387b2_fcb43823,
        64'hfca43c23_0080f822,
        64'hfc067139_80826105,
        64'h644260e2_0001e8df,
        64'hf0ef853e_85bafea4,
        64'h47039381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef40523,
        64'h87bafef4_05a387b6,
        64'hfef42623_873286ae,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e2853e_87aae7ff,
        64'hf0ef853e_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h05a387ba_fef42623,
        64'h872e87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_0001f39f,
        64'hf0ef853e_85bafe84,
        64'h57039381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef41423,
        64'h87bafef4_05a387b6,
        64'hfef42623_873286ae,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e2853e_87aaf1df,
        64'hf0ef853e_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h05a387ba_fef42623,
        64'h872e87aa_1000e822,
        64'hec061101_80826145,
        64'h74220001_c398fd44,
        64'h2703fe84_3783fef4,
        64'h3423fd84_3783fcf4,
        64'h2a2387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61457422_000100e7,
        64'h9023fd64_5703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_1b2387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61457422,
        64'h000100e7_8023fd74,
        64'h4703fe84_3783fef4,
        64'h3423fd84_3783fcf4,
        64'h0ba387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61056462_853e2781,
        64'h439cfe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826105_6462853e,
        64'h93c117c2_0007d783,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61056462_853e0ff7,
        64'hf7930007_c783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826145,
        64'h7422853e_fe843783,
        64'hfae7f5e3_47850007,
        64'h871bfe44_2783fef4,
        64'h22232785_fe442783,
        64'ha829fef4_342397ba,
        64'h1c870713_1ffee717,
        64'h078a97ba_078e87ba,
        64'hfe446703_02f71063,
        64'h27812701_fde45703,
        64'h0007d783_97ba1fa6,
        64'h8713078a_97ba078e,
        64'h87bafe44_67031ffe,
        64'he697a0b9_fe042223,
        64'hfe043423_fcf41f23,
        64'h87aa1800_f4227179,
        64'h80826145_740270a2,
        64'h0001fef7_68e3fe04,
        64'h3783fe84_3703fea4,
        64'h3423fbff_f0effef4,
        64'h302397ba_fe843783,
        64'h873e078a_97ba078a,
        64'h87bafd84_3703fea4,
        64'h3423fdff_f0effca4,
        64'h3c231800_f022f406,
        64'h71798082_01416422,
        64'h853e639c_17e10200,
        64'hc7b70800_e4221141,
        64'h80826109_640660a6,
        64'h853efec4_2783fef4,
        64'h262387aa_b38ff0ef,
        64'hc2650513_fffff517,
        64'h85be567d_fb843683,
        64'hfd040793_fe043703,
        64'hfcf43c23_fc043783,
        64'hfcf43823_fc843783,
        64'hfef43023_fd878793,
        64'h03040793_03143423,
        64'h03043023_ec1ce818,
        64'he414fac4_3c23fcb4,
        64'h3023fca4_34230880,
        64'he0a2e486_71198082,
        64'h61457402_70a2853e,
        64'h87aab9ef_f0efbf65,
        64'h0513ffff_f517fe84,
        64'h3583fe04_3603fd84,
        64'h3683fd04_3703fcd4,
        64'h3823fcc4_3c23feb4,
        64'h3023fea4_34231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'h87aabdef_f0efc945,
        64'h0513ffff_f51785be,
        64'h567dfd84_3683fd04,
        64'h3703fe84_0793fcb4,
        64'h3823fca4_3c231800,
        64'hf022f406_71798082,
        64'h61657442_70e2853e,
        64'hfec42783_fef42623,
        64'h87aac1ef_f0efc765,
        64'h0513ffff_f517fd84,
        64'h3583fd04_3603fc84,
        64'h3683873e_fe043783,
        64'hfef43023_fd878793,
        64'h03040793_03143423,
        64'h03043023_ec1ce818,
        64'he414fcc4_3423fcb4,
        64'h3823fca4_3c230080,
        64'hf822fc06_71598082,
        64'h61257402_70a2853e,
        64'hfec42783_fef42623,
        64'h87aac7ef_f0efcd65,
        64'h0513ffff_f517fd84,
        64'h3583567d_fd043683,
        64'h873efe04_3783fef4,
        64'h3023fd07_87930304,
        64'h07930314_34230304,
        64'h3023ec1c_e818e414,
        64'he010fcb4_3823fca4,
        64'h3c231800_f022f406,
        64'h711d8082_61097442,
        64'h70e2853e_fec42783,
        64'hfef42623_87aacdaf,
        64'hf0efd905_0513ffff,
        64'hf51785be_567dfc84,
        64'h3683fd84_0793fe04,
        64'h3703fef4_3023fc87,
        64'h87930404_07930314,
        64'h3c230304_3823f41c,
        64'hf018ec14_e810e40c,
        64'hfca43423_0080f822,
        64'hfc067119_8082610d,
        64'h644a60ea_853e2781,
        64'hfd843783_97024501,
        64'hf9043583_863ef884,
        64'h3683f984_3703fd84,
        64'h3783a019_17fdf884,
        64'h378300f7_6663f884,
        64'h3783fd84_3703d807,
        64'h99630007_c783f804,
        64'h37830001_f8f43023,
        64'h0785f804_37839702,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h37830007_c503f804,
        64'h3783a80d_f8f43023,
        64'h0785f804_37839702,
        64'h02500513_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_3783a8b9,
        64'hf8f43023_0785f804,
        64'h3783fca4_3c23ba2f,
        64'hf0eff984_3503f904,
        64'h3583fd84_3603f884,
        64'h36838736_47814841,
        64'h88bae03e_fe842783,
        64'he43efec4_2783fe44,
        64'h270386be_639cf6e4,
        64'h3c230087_8713f784,
        64'h3783a089_fca43c23,
        64'hcfcff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_87364781,
        64'h484188ba_e03efe84,
        64'h2783e43e_fec42783,
        64'hfe442703_86be639c,
        64'hf6e43c23_00878713,
        64'hf7843783_c3b10ff7,
        64'hf793fbb4_4783faf4,
        64'h0da34785_fef42623,
        64'h0217e793_fec42783,
        64'hfef42423_47c1a239,
        64'hf8f43023_0785f804,
        64'h3783fce7_e7e32701,
        64'hfe842703_fce42223,
        64'h0017871b_fc442783,
        64'h97020200_0513f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'ha00dcf8d_27818b89,
        64'hfec42783_fbcdfee4,
        64'h2223fff7_871bfe44,
        64'h2783d3e1_27814007,
        64'hf793fec4_2783cf91,
        64'h0007c783_fc843783,
        64'h9702f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_0007c503,
        64'hfce43423_00178713,
        64'hfc843783_a03dfce7,
        64'he7e32701_fe842703,
        64'hfce42223_0017871b,
        64'hfc442783_97020200,
        64'h0513f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_a00de7a5,
        64'h27818b89_fec42783,
        64'hfcf42223_87b200d7,
        64'h73630006_071b0007,
        64'h869bfe44_2783fc44,
        64'h2603cf91_27814007,
        64'hf793fec4_2783fcf4,
        64'h222387aa_8aaff0ef,
        64'hfc843503_85be57fd,
        64'ha011fe44_6783c781,
        64'h2781fe44_2783fcf4,
        64'h3423639c_f6e43c23,
        64'h00878713_f7843783,
        64'ha4a1f8f4_30230785,
        64'hf8043783_fce7e7e3,
        64'h2701fe84_2703fce4,
        64'h28230017_871bfd04,
        64'h27839702_02000513,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h3783a00d_cf8d2781,
        64'h8b89fec4_27839702,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h37830ff7_f513439c,
        64'hf6e43c23_00878713,
        64'hf7843783_fce7e7e3,
        64'h2701fe84_2703fce4,
        64'h28230017_871bfd04,
        64'h27839702_02000513,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h3783a00d_ef8d2781,
        64'h8b89fec4_2783fcf4,
        64'h28234785_a631f8f4,
        64'h30230785_f8043783,
        64'hfca43c23_e50ff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h47818836_88b2e03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_2603fd44,
        64'h6683fb44_6703faf4,
        64'h2a232781_439cf6e4,
        64'h3c230087_8713f784,
        64'h3783a801_278193c1,
        64'h17c2439c_f6e43c23,
        64'h00878713_f7843783,
        64'hcf812781_0807f793,
        64'hfec42783_a8152781,
        64'h0ff7f793_439cf6e4,
        64'h3c230087_8713f784,
        64'h3783cf81_27810407,
        64'hf793fec4_2783a841,
        64'hfca43c23_ee0ff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h47818836_88b2e03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_2603fd44,
        64'h66836398_f6e43c23,
        64'h00878713_f7843783,
        64'hc3b12781_1007f793,
        64'hfec42783_a8f9fca4,
        64'h3c23847f_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_36834781,
        64'h883688b2_e03efe84,
        64'h2783e43e_fec42783,
        64'hfe442603_fd446683,
        64'h6398f6e4_3c230087,
        64'h8713f784_3783c3b1,
        64'h27812007_f793fec4,
        64'h2783a235_fca43c23,
        64'hf7cff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_87b68832,
        64'h88aee03e_fe842783,
        64'he43efec4_2783fe44,
        64'h2583fd44_66030ff7,
        64'hf69301f7_d79bfb04,
        64'h27839301_02079713,
        64'h27812781_40f707bb,
        64'h8f3dfb04_270341f7,
        64'hd79bfb04_2783faf4,
        64'h2823439c_f6e43c23,
        64'h00878713_f7843783,
        64'ha8012781_4107d79b,
        64'h0107979b_439cf6e4,
        64'h3c230087_8713f784,
        64'h3783cf91_27810807,
        64'hf793fec4_2783a81d,
        64'h27810ff7_f793439c,
        64'hf6e43c23_00878713,
        64'hf7843783_cf812781,
        64'h0407f793_fec42783,
        64'ha2cdfca4_3c23833f,
        64'hf0eff984_3503f904,
        64'h3583fd84_3603f884,
        64'h3683872e_87ba8836,
        64'h88b2e03e_fe842783,
        64'he43efec4_2783fe44,
        64'h2603fd44_66830ff7,
        64'hf71393fd_fa843783,
        64'h85be8f99_8fb9fa84,
        64'h378343f7_d713fa84,
        64'h3783faf4_3423639c,
        64'hf6e43c23_00878713,
        64'hf7843783_c3bd2781,
        64'h1007f793_fec42783,
        64'hac89fca4_3c239bbf,
        64'hf0eff984_3503f904,
        64'h3583fd84_3603f884,
        64'h3683872e_87ba8836,
        64'h88b2e03e_fe842783,
        64'he43efec4_2783fe44,
        64'h2603fd44_66830ff7,
        64'hf71393fd_fa043783,
        64'h85be8f99_8fb9fa04,
        64'h378343f7_d713fa04,
        64'h3783faf4_3023639c,
        64'hf6e43c23_00878713,
        64'hf7843783_c3bd2781,
        64'h2007f793_fec42783,
        64'h18f71d63_06400793,
        64'h873e0007_c783f804,
        64'h378300f7_0b630690,
        64'h0793873e_0007c783,
        64'hf8043783_fef42623,
        64'h9bf9fec4_2783c791,
        64'h27814007_f793fec4,
        64'h2783fef4_26239bcd,
        64'hfec42783_00f70763,
        64'h06400793_873e0007,
        64'hc783f804_378302f7,
        64'h00630690_0793873e,
        64'h0007c783_f8043783,
        64'hfef42623_0207e793,
        64'hfec42783_00f71863,
        64'h05800793_873e0007,
        64'hc783f804_3783fef4,
        64'h26239bbd_fec42783,
        64'hfcf42a23_47a9a809,
        64'hfcf42a23_478900f7,
        64'h16630620_0793873e,
        64'h0007c783_f8043783,
        64'ha035fcf4_2a2347a1,
        64'h00f71663_06f00793,
        64'h873e0007_c783f804,
        64'h3783a099_fcf42a23,
        64'h47c100f7_16630580,
        64'h0793873e_0007c783,
        64'hf8043783_00f70b63,
        64'h07800793_873e0007,
        64'hc783f804_37838782,
        64'h97bac1a7_87930000,
        64'h57970007_871b439c,
        64'h97bac2a7_87930000,
        64'h57970027_97139381,
        64'h02069793_6ce7e363,
        64'h05300793_0006871b,
        64'hfdb7869b_27810007,
        64'hc783f804_37830001,
        64'ha0110001_a0210001,
        64'ha031f8f4_30230785,
        64'hf8043783_fef42623,
        64'h1007e793_fec42783,
        64'ha015f8f4_30230785,
        64'hf8043783_fef42623,
        64'h1007e793_fec42783,
        64'ha835f8f4_30230785,
        64'hf8043783_fef42623,
        64'h1007e793_fec42783,
        64'ha889f8f4_30230785,
        64'hf8043783_fef42623,
        64'h0407e793_fec42783,
        64'h06f71663_06800793,
        64'h873e0007_c783f804,
        64'h3783f8f4_30230785,
        64'hf8043783_fef42623,
        64'h0807e793_fec42783,
        64'ha079f8f4_30230785,
        64'hf8043783_fef42623,
        64'h2007e793_fec42783,
        64'h0af71463_06c00793,
        64'h873e0007_c783f804,
        64'h3783f8f4_30230785,
        64'hf8043783_fef42623,
        64'h1007e793_fec42783,
        64'h878297ba_ce078793,
        64'h00005797_0007871b,
        64'h439c97ba_cf078793,
        64'h00005797_00279713,
        64'h93810206_97930ee7,
        64'he96347c9_0006871b,
        64'hf987869b_27810007,
        64'hc783f804_3783f8f4,
        64'h30230785_f8043783,
        64'hfef42223_27814781,
        64'h00075363_0007871b,
        64'hfbc42783_faf42e23,
        64'h439cf6e4_3c230087,
        64'h8713f784_378302f7,
        64'h1a6302a0_0793873e,
        64'h0007c783_f8043783,
        64'ha091fef4_222387aa,
        64'hf86ff0ef_853ef804,
        64'h0793cb91_87aaf54f,
        64'hf0ef853e_0007c783,
        64'hf8043783_f8f43023,
        64'h0785f804_3783fef4,
        64'h26234007_e793fec4,
        64'h278308f7_106302e0,
        64'h0793873e_0007c783,
        64'hf8043783_fe042223,
        64'hf8f43023_0785f804,
        64'h3783fef4_2423fc04,
        64'h2783a029_fef42423,
        64'h278140f0_07bbfc04,
        64'h2783fef4_26230027,
        64'he793fec4_27830207,
        64'hd0632781_fc042783,
        64'hfcf42023_439cf6e4,
        64'h3c230087_8713f784,
        64'h378304f7_176302a0,
        64'h0793873e_0007c783,
        64'hf8043783_a8b9fef4,
        64'h242387aa_833ff0ef,
        64'h853ef804_0793cb91,
        64'h87aa801f_f0ef853e,
        64'h0007c783_f8043783,
        64'hfe042423_f3852781,
        64'hfe042783_0001fe04,
        64'h2023a021_fef42023,
        64'h4785f8f4_30230785,
        64'hf8043783_fef42623,
        64'h0107e793_fec42783,
        64'ha01dfef4_20234785,
        64'hf8f43023_0785f804,
        64'h3783fef4_26230087,
        64'he793fec4_2783a091,
        64'hfef42023_4785f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0047e793,
        64'hfec42783_a08dfef4,
        64'h20234785_f8f43023,
        64'h0785f804_3783fef4,
        64'h26230027_e793fec4,
        64'h2783a041_fef42023,
        64'h4785f8f4_30230785,
        64'hf8043783_fef42623,
        64'h0017e793_fec42783,
        64'h878297ba_e9478793,
        64'h00005797_0007871b,
        64'h439c97ba_ea478793,
        64'h00005797_00279713,
        64'h93810206_97930ce7,
        64'he06347c1_0006871b,
        64'hfe07869b_27810007,
        64'hc783f804_3783fe04,
        64'h2623f8f4_30230785,
        64'hf8043783_2270006f,
        64'hf8f43023_0785f804,
        64'h37839702_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_37830007,
        64'hc503f804_378302f7,
        64'h0b630250_0793873e,
        64'h0007c783_f8043783,
        64'h26b0006f_f8f43c23,
        64'h86678793_00000797,
        64'h26079de3_f9043783,
        64'hfc043c23_f6e43c23,
        64'hf8d43023_f8c43423,
        64'hf8b43823_f8a43c23,
        64'h1100e922_ed067135,
        64'h8082610d_644a60ea,
        64'h853e87aa_b47ff0ef,
        64'hfb843503_fb043583,
        64'hfa843603_fa043683,
        64'hfe843783_883688b2,
        64'he03ef904_2783e43e,
        64'h401ce83e_441cfc04,
        64'h0713f974_46830007,
        64'h861bf884_3783f6e7,
        64'hffe347fd_fe843703,
        64'hc791f984_3783f8f4,
        64'h3c2302f7_57b3f884,
        64'h3783f984_3703fcf7,
        64'h08239736_ff040693,
        64'hfed43423_00170693,
        64'hfe843703_0ff7f793,
        64'h37d90ff7_f7939fb9,
        64'hfe744703_06100793,
        64'ha0190410_0793c781,
        64'h27810207_f793441c,
        64'ha01d0ff7_f7930307,
        64'h879bfe74_478300e7,
        64'he96347a5_0ff7f713,
        64'hfe744783_fef403a3,
        64'h02f777b3_f8843783,
        64'hf9843703_c7c1f984,
        64'h3783c781_27814007,
        64'hf793441c_c41c9bbd,
        64'h441ce781_f9843783,
        64'hfe043423_f8f42823,
        64'h87baf8f4_0ba38746,
        64'hf9043423_f8e43c23,
        64'hfad43023_fac43423,
        64'hfab43823_faa43c23,
        64'h1100e922_ed067135,
        64'h8082610d_644a60ea,
        64'h853e87aa_c5fff0ef,
        64'hfb843503_fb043583,
        64'hfa843603_fa043683,
        64'hfe843783_883688b2,
        64'he03ef904_2783e43e,
        64'h401ce83e_441cfc04,
        64'h0713f974_46830007,
        64'h861bf884_3783f6e7,
        64'hffe347fd_fe843703,
        64'hc791f984_3783f8f4,
        64'h3c2302f7_57b3f884,
        64'h3783f984_3703fcf7,
        64'h08239736_ff040693,
        64'hfed43423_00170693,
        64'hfe843703_0ff7f793,
        64'h37d90ff7_f7939fb9,
        64'hfe744703_06100793,
        64'ha0190410_0793c781,
        64'h27810207_f793441c,
        64'ha01d0ff7_f7930307,
        64'h879bfe74_478300e7,
        64'he96347a5_0ff7f713,
        64'hfe744783_fef403a3,
        64'h02f777b3_f8843783,
        64'hf9843703_c7c1f984,
        64'h3783c781_27814007,
        64'hf793441c_c41c9bbd,
        64'h441ce781_f9843783,
        64'hfe043423_f8f42823,
        64'h87baf8f4_0ba38746,
        64'hf9043423_f8e43c23,
        64'hfad43023_fac43423,
        64'hfab43823_faa43c23,
        64'h1100e922_ed067135,
        64'h80826161_640660a6,
        64'h853e87aa_c65ff0ef,
        64'hfe843503_fe043583,
        64'hfd843603_fd043683,
        64'hfc843703_fc043783,
        64'h883e88ba_441c4818,
        64'h00e78023_02000713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h3783cf91_27818ba1,
        64'h481ca015_00e78023,
        64'h02b00713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_3783cf99,
        64'h27818b91_481ca0a1,
        64'h00e78023_02d00713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h3783cf99_0ff7f793,
        64'hfbf44783_06e7e863,
        64'h47fdfc04_370300e7,
        64'h80230300_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'h00e7ef63_47fdfc04,
        64'h370300e7_80230620,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_00e7ef63,
        64'h47fdfc04_370302f7,
        64'h14634789_0007871b,
        64'hfb842783_a81500e7,
        64'h80230580_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'h02e7e063_47fdfc04,
        64'h3703c785_27810207,
        64'hf793481c_02f71a63,
        64'h47c10007_871bfb84,
        64'h2783a88d_00e78023,
        64'h07800713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_378302e7,
        64'he06347fd_fc043703,
        64'he7852781_0207f793,
        64'h481c02f7_1a6347c1,
        64'h0007871b_fb842783,
        64'hfcf43023_17fdfc04,
        64'h378300f7_176347c1,
        64'h0007871b_fb842783,
        64'hcf89fc04_3783fcf4,
        64'h302317fd_fc043783,
        64'h02f71663_fc043703,
        64'h00846783_00f70863,
        64'hfc043703_00046783,
        64'hc3a9fc04_3783e7a1,
        64'h27814007_f793481c,
        64'h12078363_27818bc1,
        64'h481cfce7_f6e347fd,
        64'hfc043703_00f77763,
        64'hfc043703_00846783,
        64'hcf812781_8b85481c,
        64'h00e78023_03000713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h3783a831_fce7fae3,
        64'h47fdfc04_370302f7,
        64'h7563fc04_37030004,
        64'h678300e7_80230300,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_a831c41c,
        64'h37fd441c_c3952781,
        64'h8bb1481c_e7890ff7,
        64'hf793fbf4_4783cb9d,
        64'h27818b85_481ccf9d,
        64'h2781441c_ebd12781,
        64'h8b89481c_faf42c23,
        64'h87bafaf4_0fa38746,
        64'h87c2fcf4_3023fce4,
        64'h3423fcd4_3823fcc4,
        64'h3c23feb4_3023fea4,
        64'h34230880_e0a2e486,
        64'h715d8082_61256446,
        64'h60e6853e_fc843783,
        64'hfcf769e3_fac46783,
        64'h8f1dfe04_3783fc84,
        64'h37039702_02000513,
        64'hfd043583_863efc04,
        64'h3683fd84_3703fce4,
        64'h34230017_8713fc84,
        64'h3783a00d_cb9d2781,
        64'h8b89fa84_2783f7e1,
        64'hfb043783_9702fd04,
        64'h3583863e_fc043683,
        64'hfd843703_fce43423,
        64'h00178713_fc843783,
        64'h0007c503_97bafb04,
        64'h3783fb84_3703faf4,
        64'h382317fd_fb043783,
        64'ha81dfcf7_67e3fe84,
        64'h3703fac4_6783fef4,
        64'h34230785_fe843783,
        64'h97020200_0513fd04,
        64'h3583863e_fc043683,
        64'hfd843703_fce43423,
        64'h00178713_fc843783,
        64'ha035fef4_3423fb04,
        64'h3783efa5_27818b85,
        64'hfa842783_e3c92781,
        64'h8b89fa84_2783fef4,
        64'h3023fc84_3783faf4,
        64'h242387ba_faf42623,
        64'h874687c2_faf43823,
        64'hfae43c23_fcd43023,
        64'hfcc43423_fcb43823,
        64'hfca43c23_1080e8a2,
        64'hec86711d_80826145,
        64'h740270a2_853efec4,
        64'h2783ffc5_87aaf6df,
        64'hf0ef853e_0007c783,
        64'h639cfd84_3783fef4,
        64'h2623fd07_879b2781,
        64'h9fb92781_0007c783,
        64'he290fd84_36830017,
        64'h8613639c_fd843783,
        64'h0007871b_0017979b,
        64'h9fb90027_979b87ba,
        64'hfec42703_a825fe04,
        64'h2623fca4_3c231800,
        64'hf022f406_71798082,
        64'h61056462_853e0ff7,
        64'hf7938b85_4781a011,
        64'h478500e7_e4630390,
        64'h07930ff7_f713fef4,
        64'h478300e7_fc6302f0,
        64'h07930ff7_f713fef4,
        64'h4783fef4_07a387aa,
        64'h1000ec22_11018082,
        64'h61457422_853e2781,
        64'h40f707b3_fd843783,
        64'hfe843703_f3e5fce4,
        64'h3823fff7_8713fd04,
        64'h3783cb81_0007c783,
        64'hfe843783_fef43423,
        64'h0785fe84_3783a031,
        64'hfef43423_fd843783,
        64'hfcb43823_fca43c23,
        64'h1800f422_71798082,
        64'h61457402_70a20001,
        64'h9682853e_85bafef4,
        64'h47836798_fe043783,
        64'h6394fe04_3783cf81,
        64'h0ff7f793_fef44783,
        64'hfef407a3_fcd43823,
        64'hfcc43c23_feb43023,
        64'h87aa1800_f022f406,
        64'h71798082_61457402,
        64'h70a20001_8e7ff0ef,
        64'h853efef4_4783c791,
        64'h0ff7f793_fef44783,
        64'hfef407a3_fcd43823,
        64'hfcc43c23_feb43023,
        64'h87aa1800_f022f406,
        64'h71798082_61457422,
        64'h0001fef4_07a3fcd4,
        64'h3823fcc4_3c23feb4,
        64'h302387aa_1800f422,
        64'h71798082_61457422,
        64'h000100e7_8023fef4,
        64'h470397ba_fd843783,
        64'hfe043703_00f77b63,
        64'hfd043783_fd843703,
        64'hfef407a3_fcd43823,
        64'hfcc43c23_feb43023,
        64'h87aa1800_f4227179,
        64'h8082610d_690a64aa,
        64'h644a60ea_f6040113,
        64'h853e8126_814a4781,
        64'h2b0010ef_71c50513,
        64'h00005517_a80157f9,
        64'h2c0010ef_4dc50513,
        64'h00005517_85befac4,
        64'h27832d20_10ef4d65,
        64'h05130000_5517c395,
        64'h2781fac4_2783faf4,
        64'h262387aa_b63ff0ef,
        64'hf6843503_85be863a,
        64'hf6442703_2781739c,
        64'hf8043783_304010ef,
        64'h75850513_00005517,
        64'hf8f43023_f8843783,
        64'heae7d2e3_478d0007,
        64'h871bfd04_2783fcf4,
        64'h28232785_fd042783,
        64'h330010ef_5a450513,
        64'h00005517_fce7d6e3,
        64'h04700793_0007871b,
        64'hfdc42783_fcf42e23,
        64'h2785fdc4_27833560,
        64'h10ef7225_05130000,
        64'h551785be_27810387,
        64'hc78397ba_fdc42783,
        64'hf7843703_a02dfc04,
        64'h2e2337a0_10ef7b65,
        64'h05130000_55173860,
        64'h10ef7aa5_05130000,
        64'h551785be_7b9cf784,
        64'h378339a0_10ef7a65,
        64'h05130000_551785be,
        64'h779cf784_37833ae0,
        64'h10ef7a25_05130000,
        64'h551785be_739cf784,
        64'h3783fce7_d7e347bd,
        64'h0007871b_fd842783,
        64'hfcf42c23_2785fd84,
        64'h27833da0_10ef7a65,
        64'h05130000_551785be,
        64'h27810107_c78397ba,
        64'hfd842783_f7843703,
        64'ha02dfc04_2c233fe0,
        64'h10ef7d25_05130000,
        64'h5517fce7_d7e347bd,
        64'h0007871b_fd442783,
        64'hfcf42a23_2785fd44,
        64'h27834220_10ef7ee5,
        64'h05130000_551785be,
        64'h27810007_c78397ba,
        64'hfd442783_f7843703,
        64'ha02dfc04_2a234460,
        64'h10ef7f25_05130000,
        64'h55174520_10ef7e65,
        64'h05130000_551785be,
        64'hfd042783_f6f43c23,
        64'h97ba2701_0077171b,
        64'hfd042703_f8843783,
        64'haa91fc04_2823aac9,
        64'h57f94820_10ef7f65,
        64'h05130000_551785be,
        64'hfac42783_494010ef,
        64'h69850513_00005517,
        64'hc3952781_fac42783,
        64'hfaf42623_87aad25f,
        64'hf0ef853a_85be4605,
        64'h278167bc_fa043783,
        64'hf8843703_f8f43423,
        64'h00078793_878a40f1,
        64'h01330792_839107bd,
        64'hf8e43823_177d873e,
        64'h893a870a_fc043783,
        64'h4e8010ef_83c50513,
        64'h00006517_85be4bfc,
        64'hfa043783_4fc010ef,
        64'h83050513_00006517,
        64'h85be4bbc_fa043783,
        64'h510010ef_81c50513,
        64'h00006517_85be67bc,
        64'hfa043783_524010ef,
        64'h81850513_00006517,
        64'h85be739c_fa043783,
        64'h538010ef_81450513,
        64'h00006517_85be6f9c,
        64'hfa043783_54c010ef,
        64'h81050513_00006517,
        64'h85be4bdc_fa043783,
        64'h560010ef_80c50513,
        64'h00006517_85be4b9c,
        64'hfa043783_574010ef,
        64'h80850513_00006517,
        64'h85be47dc_fa043783,
        64'h588010ef_80450513,
        64'h00006517_85be479c,
        64'hfa043783_59c010ef,
        64'h81050513_00006517,
        64'hfce7d7e3_479d0007,
        64'h871bfcc4_2783fcf4,
        64'h26232785_fcc42783,
        64'h5c0010ef_82c50513,
        64'h00006517_85be2781,
        64'h0007c783_97baf984,
        64'h3703fcc4_2783a02d,
        64'hfc042623_f8f43c23,
        64'hfa043783_5ec010ef,
        64'h84850513_00006517,
        64'h5f8010ef_83450513,
        64'h00006517_faf43023,
        64'hfb043783_a68d57f9,
        64'h610010ef_82c50513,
        64'h00006517_85befac4,
        64'h27836220_10ef8265,
        64'h05130000_6517c395,
        64'h2781fac4_2783faf4,
        64'h262387aa_eb3ff0ef,
        64'h853e4585_4605fb04,
        64'h3783faf4_38230007,
        64'h8793878a_40f10133,
        64'h07928391_07bdfae4,
        64'h3c23177d_873efc04,
        64'h3783fcf4_30232000,
        64'h07936720_10ef85e5,
        64'h05130000_6517aed1,
        64'h57fd6820_10ef8465,
        64'h05130000_6517cb89,
        64'h2781fc84_2783fcf4,
        64'h242387aa_e5bff0ef,
        64'h84be878a_f6f42223,
        64'h87aef6a4_34231100,
        64'he14ae526_e922ed06,
        64'h71358082_61457402,
        64'h70a2853e_4781a011,
        64'h57fd6ca0_10ef86e5,
        64'h05130000_651785be,
        64'hfe442783_cf812781,
        64'hfe442783_fef42223,
        64'h87aa7600_30efc5e5,
        64'h05131fff_051785be,
        64'h863afe84_3683fd44,
        64'h2783fd04_2703fae7,
        64'he0e3678d_0007871b,
        64'hfd042783_fef43423,
        64'h97ba0060_07b7fe84,
        64'h3703fcf4_28239fb9,
        64'h77f5fd04_2703a0b5,
        64'h57fd7320_10ef8d65,
        64'h05130000_651785be,
        64'hfe042783_cf812781,
        64'hfe042783_fef42023,
        64'h87aa7c80_30efcc65,
        64'h05131fff_051785be,
        64'h660dfe84_3683fd44,
        64'h2783a8a1_fef43423,
        64'hfd843783_fcf42823,
        64'h87bafcf4_2a238732,
        64'h87aefca4_3c231800,
        64'hf022f406_71798082,
        64'h61056442_60e2853e,
        64'h478179a0_10ef91e5,
        64'h05130000_6517a801,
        64'h57f57aa0_10ef8fe5,
        64'h05130000_651785be,
        64'hfe442783_cf812781,
        64'hfe442783_fef42223,
        64'h87aa53c0_20efd3e5,
        64'h05131fff_0517a081,
        64'h57f97da0_10ef9065,
        64'h05130000_651785be,
        64'hfe442783_cf812781,
        64'hfe442783_fef42223,
        64'h87aa4ab0_10efd6e5,
        64'h05131fff_0517fe84,
        64'h3583863e_43dcfe84,
        64'h3783a8b5_57fd0170,
        64'h10ef9225_05130000,
        64'h6517eb89_fe843783,
        64'hfea43423_289010ef,
        64'h45010330_10ef9265,
        64'h05130000_65171000,
        64'he822ec06_11018082,
        64'h61457402_70a20001,
        64'heb9ff0ef_01078513,
        64'h07fa478d_02000593,
        64'hec9ff0ef_00878513,
        64'h07fa478d_0c700593,
        64'hed9ff0ef_00c78513,
        64'h07fa478d_458dee7f,
        64'hf0ef0047_851307fa,
        64'h478d85be_0ff7f793,
        64'h27810087_d79bfec4,
        64'h2783f03f_f0ef01e7,
        64'h9513478d_85be0ff7,
        64'hf793fec4_2783f17f,
        64'hf0ef00c7_851307fa,
        64'h478d0800_0593f27f,
        64'hf0ef0047_851307fa,
        64'h478d4581_fef42623,
        64'h02f757bb_fdc42703,
        64'h27810047_979bfd84,
        64'h2783fcf4_2c2387ba,
        64'hfcf42e23_872e87aa,
        64'h1800f022_f4067179,
        64'h80826105_644260e2,
        64'h0001f6bf_f0ef01e7,
        64'h9513478d_85befef4,
        64'h4783dfed_87aafc9f,
        64'hf0ef0001_fef407a3,
        64'h87aa1000_e822ec06,
        64'h11018082_01416402,
        64'h60a2853e_27810207,
        64'hf7932781_87aafd3f,
        64'hf0ef0147_851307fa,
        64'h478d0800_e022e406,
        64'h11418082_61056462,
        64'h853e0ff7_f7930007,
        64'hc783fe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826145_74220001,
        64'h00e78023_fd744703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf40ba3,
        64'h87aefca4_3c231800,
        64'hf4227179_a00119f0,
        64'h10efa6a5_05130000,
        64'h65178402_03c58593,
        64'h00006597_10000437,
        64'heb812781_fe442783,
        64'h1c1010ef_a6450513,
        64'h00006517_fce7d7e3,
        64'h47bd0007_871bfe84,
        64'h2783fef4_24232785,
        64'hfe842783_1e5010ef,
        64'haa850513_00006517,
        64'h85be2781_0007c783,
        64'h97bafd84_3703fe84,
        64'h2783a02d_fe042423,
        64'h209010ef_ab450513,
        64'h00006517_100005b7,
        64'hfcf43c23_100007b7,
        64'hfef42223_87aa3700,
        64'h00ef1000_053765a1,
        64'h231010ef_ad450513,
        64'h00006517_fce7dae3,
        64'h47890007_871bfec4,
        64'h2783fef4_26232785,
        64'hfec42783_255010ef,
        64'haf050513_00006517,
        64'h473010ef_24078513,
        64'h000f47b7_a015fe04,
        64'h26232730_10efae65,
        64'h05130000_651718a0,
        64'h00efa007_85130262,
        64'h67b72007_859367f1,
        64'h1800f022_f4067179,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_100004b7,
        64'h15058593_00006597,
        64'hf1402573_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_090000ef,
        64'hf9810113_3fff0117,
        64'hfeb56ce3_00450513,
        64'h00052023_00b57863,
        64'hc4218593_ffc50513,
        64'h1fff0517_fec5e8e3,
        64'h00458593_00450513,
        64'h0055a023_00052283,
        64'h00c5fc63_01c60613,
        64'h1fff0617_fdc58593,
        64'h1fff0597_de450513,
        64'h00007517_83418193,
        64'h1fff1197_09249063,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
