/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 2098;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00000078_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000078_36313025,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000078_36313025,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_78323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000a64_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h00000a64_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_0000000a,
        64'h78363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h0000000a_78363130,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h0000000a_78363130,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_00000a64,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_00000a64,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_00000a64,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_00000a64,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h00000000_00000a78,
        64'h25202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h00000000_0000000a,
        64'h2164656c_69616620,
        64'h64616552_20304453,
        64'h0000000a_21206465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_0a212064,
        64'h656c6961_66206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a2120,
        64'h64656c69_61662067,
        64'h69666e6f_43204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_002e2e2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd0080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h08090000_38000000,
        64'hda0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000a001,
        64'h830fe0ef_1bc50513,
        64'h00001517_84025b65,
        64'h85930000_05971000,
        64'h0437e901_dcafd0ef,
        64'h10000537_65a1856f,
        64'he0ef1da5_05130000,
        64'h1517950f_e0ef2404,
        64'h051386af_e0ef1ee5,
        64'h05130000_1517964f,
        64'he0ef2404_0513000f,
        64'h4437882f_e0ef1de5,
        64'h05130000_1517d30f,
        64'hd0efe022_e406a005,
        64'h05132005_85931141,
        64'h02626537_65f18082,
        64'h0141421c_920100f6,
        64'h90231602_47892641,
        64'h640260a2_80820141,
        64'h45056402_60a28082,
        64'h01414505_00f61023,
        64'h3ff7879b_920177fd,
        64'h16026402_60a20326,
        64'h061bfe07_56e38b89,
        64'h4107571b_0107971b,
        64'h93c117c2_0006d783,
        64'hef9da011_92811682,
        64'h0306069b_4050e129,
        64'hde0fe0ef_842ae406,
        64'he0226000_05934681,
        64'h862e1141_80820141,
        64'h439c9381_00e69023,
        64'h17824709_0106079b,
        64'h640260a2_80820141,
        64'h450562e7_ac234705,
        64'h00000797_640260a2,
        64'h948fe0ef_63c50513,
        64'h65058593_35c00613,
        64'h00001517_00001597,
        64'h80820141_45056402,
        64'h60a28082_01414505,
        64'h66e7a723_47050000,
        64'h07976402_60a297ef,
        64'he0ef6725_05136865,
        64'h859335d0_06130000,
        64'h15170000_15978082,
        64'h01414505_00e79023,
        64'h3ff7071b_9381777d,
        64'h17826402_60a20326,
        64'h079bfe07_56e38b89,
        64'h4107571b_0107971b,
        64'h93c117c2_0006d783,
        64'hebd9a011_92811682,
        64'h0306069b_4050e53d,
        64'heb0fe0ef_6ee79423,
        64'h85228005_85934601,
        64'h46854745_00000797,
        64'h6585c0df_e0ef8522,
        64'h458500e7_90239381,
        64'h17822791_862e2000,
        64'h0713405c_fee79de3,
        64'h07850007_802308d6,
        64'h12632005_871387ae,
        64'h842a1116_86937207,
        64'ha3231111_16b70000,
        64'h07975150_c979e022,
        64'he4061141_80820141,
        64'h853e4785_74e7a123,
        64'h47050000_07976402,
        64'h60a2a52f_e0ef7465,
        64'h051375a5_859332c0,
        64'h06130000_15170000,
        64'h15978082_0141853e,
        64'h00a037b3_640260a2,
        64'hf50fe0ef_a0058593,
        64'h46014681_852265ad,
        64'hf17d4785_f64fe0ef,
        64'h70058593_4681658d,
        64'h49308082_0141853e,
        64'h640260a2_47857ae7,
        64'ha2234705_00000797,
        64'hab0fe0ef_7a450513,
        64'h7b858593_32d00613,
        64'h00001517_00001597,
        64'h02f70963_842a1117,
        64'h87931111_17b77c07,
        64'haa235158_00000797,
        64'hcd25e022_e4061141,
        64'hbd85bd8f_e0ef4505,
        64'hdc0780e3_0807f793,
        64'h0007d783_b3f14505,
        64'h7ee7af23_47050000,
        64'h0797b0af_e0ef7fe5,
        64'h05138125_859348e0,
        64'h06130000_15170000,
        64'h2597b7e9_ffcfe0ef,
        64'h85d2fd37_98e38522,
        64'h85ca4601_46850344,
        64'h4783c0a1_c3290407,
        64'h77130007_d7039381,
        64'h178203e7_879b405c,
        64'he20510e3_0ff4f493,
        64'h34fd833f_e0efa01d,
        64'h300a0a13_4985c54f,
        64'he0ef00e7_90230407,
        64'h67130280_0493500a,
        64'h09130007_d7039381,
        64'h88d71123_46c10000,
        64'h17171782_00d71023,
        64'h03e7879b_93011702,
        64'h0047871b_45056a05,
        64'h405c0400_069300f7,
        64'h04630800_0693478d,
        64'h03744703_08f71b63,
        64'h11178793_111117b7,
        64'h8a07af23_50580000,
        64'h1797bd69_4505d939,
        64'hc63ff0ef_85225005,
        64'h8593dc1c_031975b7,
        64'h5007879b_031977b7,
        64'h00f69023_4789bd7d,
        64'h4505dd2d_c87ff0ef,
        64'h85220805_8593dc1c,
        64'h02faf5b7_0807879b,
        64'h02faf7b7_00f69023,
        64'h4789b5a5_fe0756e3,
        64'h8b894107_571b0107,
        64'h971b93c1_17c20006,
        64'hd783ef9d_a0119281,
        64'h16820306_069b4050,
        64'hf00514e3_915fe0ef,
        64'h60000593_10060613,
        64'h468103b9_0637b5f5,
        64'h439c9381_178227c1,
        64'h405c00e7_80230047,
        64'h67130007_c7039381,
        64'h17820287_879b4501,
        64'h405cd60f_e0ef3e80,
        64'h05130af7_0a63479d,
        64'h5478f921_d17ff0ef,
        64'h852200f6_90234789,
        64'h5c0cb5e5_fe0756e3,
        64'h8b894107_571b0107,
        64'h971b93c1_17c20006,
        64'hd783efc9_a0119281,
        64'h16820306_069b4050,
        64'hf159993f_e0ef9ce7,
        64'h95238522_60000593,
        64'h16454685_47450000,
        64'h17978100_0637ef1f,
        64'he0ef4585_00e79023,
        64'h93811782_2791860a,
        64'h04000713_415c8082,
        64'h61654505_6a0669a6,
        64'h694664e6_9ee7ad23,
        64'h47050000_17977406,
        64'h70a6d0af_e0ef9fe5,
        64'h0513a125_85931f30,
        64'h06130000_25170000,
        64'h25978082_61656a06,
        64'h69a66946_64e67406,
        64'h70a64505_d135a0ff,
        64'he0ef8522_60000593,
        64'h46812006_0613dd1c,
        64'h03b90637_2007879b,
        64'h0bebc7b7_80826165,
        64'h6a0669a6_694664e6,
        64'h740670a6_4505a6e7,
        64'ha2234705_00001797,
        64'hd70fe0ef_a6450513,
        64'ha7858593_1f400613,
        64'h00002517_00002597,
        64'h80826165_45056a06,
        64'h69a66946_64e600f6,
        64'h10233ff7_879b9201,
        64'h77fd1602_740670a6,
        64'h0326061b_fe0755e3,
        64'h8b894107_571b0107,
        64'h971b93c1_17c20006,
        64'hd7831207_9a63a019,
        64'h92811682_0306069b,
        64'h4050e145_aadfe0ef,
        64'h85226000_05934681,
        64'h10060613_dd1c03b9,
        64'h06375007_879b0319,
        64'h77b70af7_0163479d,
        64'h55781ae7_88634709,
        64'h10e78b63_47050345,
        64'h478308f7_1363842a,
        64'h11178793_111117b7,
        64'hb007ab23_51580000,
        64'h17971005_0263fc02,
        64'hf802f402_f002ec02,
        64'he802e402_e002e0d2,
        64'he4cee8ca_eca6f0a2,
        64'hf4867159_80820141,
        64'h4505b4e7_a4234705,
        64'h00001797_60a2e56f,
        64'he0efb4a5_0513b5e5,
        64'h85932b70_06130000,
        64'h25170000_2597b75d,
        64'h00c69023_92411642,
        64'h8e5d0622_8fd90017,
        64'he7938205_03f7f793,
        64'h071a0096_57130006,
        64'hd783fee5_e8e32785,
        64'h92410307_961302f8,
        64'h573bf8a7_8be3a019,
        64'h7ff00513_47858082,
        64'h014100f6_90230047,
        64'he7934501_60a20006,
        64'hd783dfed_8b890006,
        64'hd78300e6_90239341,
        64'h17428f5d_0017e793,
        64'h0ff7f793_07228305,
        64'h0006d783_bfd9bee7,
        64'ha2234705_00001797,
        64'hef0fe0ef_be450513,
        64'hbf858593_2b800613,
        64'h00002517_00002597,
        64'h80820141_450560a2,
        64'hf6759341_03051713,
        64'h02f5fc63_367d0017,
        64'h151b02e8_57bb0717,
        64'h8e630365_478300f6,
        64'h902393c1_17c29be9,
        64'h93c117c2_47054625,
        64'h0006d783_92811682,
        64'h02c6869b_48890085,
        64'h28034154_04f71863,
        64'h11178793_111117b7,
        64'hc407af23_51580000,
        64'h17971005_0063e406,
        64'h11418082_0141439c,
        64'h938100e6_90231782,
        64'h47090106_079b6402,
        64'h60a28082_01414505,
        64'hc8e7a723_47050000,
        64'h17976402_60a2f9ef,
        64'he0efc925_0513ca65,
        64'h859319f0_06130000,
        64'h25170000_25978082,
        64'h01414505_640260a2,
        64'h80820141_4505cce7,
        64'ha2234705_00001797,
        64'h640260a2_fd4fe0ef,
        64'hcc850513_cdc58593,
        64'h1a000613_00002517,
        64'h00002597_80820141,
        64'h450500e7_90233ff7,
        64'h071b9381_777d1782,
        64'h640260a2_0326079b,
        64'hfe0756e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d783ebd9,
        64'ha0119281_16820306,
        64'h069b4050_e53dd07f,
        64'he0efd2e7_9f238522,
        64'h60000593_16414685,
        64'h47450000_17970100,
        64'h0637a64f_f0ef8522,
        64'h458500e7_90239381,
        64'h17822791_862e0400,
        64'h0713405c_fee79de3,
        64'h07850007_802308d6,
        64'h13630405_871387ae,
        64'h842a1116_8693d607,
        64'haf231111_16b70000,
        64'h17975150_cd61e022,
        64'he4061141_b76500e6,
        64'h90230047_67139b61,
        64'h93411742_0006d703,
        64'h92811682_03e7869b,
        64'h405cb5fd_4505d551,
        64'hd91fe0ef_85226005,
        64'h85934609_468102f4,
        64'h0ba365a1_4789f005,
        64'h15e3dabf_e0ef8522,
        64'h70058593_4681658d,
        64'h4830b7a9_4501439c,
        64'h93811782_27c1405c,
        64'h04f70163_47915478,
        64'h00e78023_0ff77713,
        64'h0206e713_00c59463,
        64'h0026e713_0ff6f693,
        64'h0007c683_93811782,
        64'h0287879b_460d0374,
        64'h4583405c_a13fe0ef,
        64'h3e800513_00f69023,
        64'h4789b725_60078613,
        64'hf2e698e3_20078613,
        64'h471102e4_0ba303b7,
        64'h07b7470d_f2f718e3,
        64'h47a14858_80820141,
        64'h4505e4e7_ac234705,
        64'h00001797_640260a2,
        64'h969fe0ef_e5c50513,
        64'he7058593_11200613,
        64'h00002517_00002597,
        64'hb7e5f4e7_e1e34501,
        64'h478d4958_b7495007,
        64'h86138082_01416402,
        64'h60a24505_e8e7ad23,
        64'h47050000_17979a7f,
        64'he0efe9a5_0513eae5,
        64'h85931130_06130000,
        64'h25170000_25978082,
        64'h01416402_60a24505,
        64'h00f61023_3ff7879b,
        64'h920177fd_16020326,
        64'h061bfe07_56e38b89,
        64'h4107571b_0107971b,
        64'h93c117c2_0006d783,
        64'he3e1a011_92811682,
        64'h0306069b_4050ed05,
        64'hed9fe0ef_85226000,
        64'h05934681_06e68f63,
        64'h10078613_471102e4,
        64'h0ba303b7_07b74709,
        64'h0ce78863_54740752,
        64'h20005737_8ff91782,
        64'h0ff78793_00ff07b7,
        64'h781814f7_0e634785,
        64'h03444703_0af70e63,
        64'h47890365_470308f7,
        64'h1a63842a_11178793,
        64'h111117b7_f407ad23,
        64'h51580000_1797c565,
        64'he022e406_1141b7a9,
        64'h439c9381_00e69023,
        64'h17824709_0106079b,
        64'h80826105_450564a2,
        64'hf8e7a323_47050000,
        64'h17976442_60e2a97f,
        64'he0eff8a5_0513f9e5,
        64'h85930b90_06130000,
        64'h25170000_2597bfb1,
        64'h450500e7_90233ff7,
        64'h071b9381_777d1782,
        64'h0326079b_fe0756e3,
        64'h8b894107_571b0107,
        64'h971b93c1_17c20006,
        64'hd783efb1_a0119281,
        64'h16820306_069b4050,
        64'hf951fc3f_e0effee7,
        64'h9d238522_30058593,
        64'h46014685_47450000,
        64'h179765ad_d1eff0ef,
        64'h85224585_00e79023,
        64'h93811782_27918626,
        64'h4721405c_80826105,
        64'h64a26442_60e24505,
        64'h02e7a323_47050000,
        64'h1797b33f_e0ef0265,
        64'h051303a5_85930ba0,
        64'h06130000_25170000,
        64'h25978082_610564a2,
        64'h644260e2_4505cd15,
        64'h830ff0ef_85227005,
        64'h85934681_658d4830,
        64'hfee79de3_07850007,
        64'h802302d6_16630085,
        64'h871387ae_84ae842a,
        64'h11168693_0807a223,
        64'h111116b7_00001797,
        64'h5150c17d_e426e822,
        64'hec061101_80826105,
        64'h450564a2_0ae7a123,
        64'h47050000_17976442,
        64'h60e2bb3f_e0ef0a65,
        64'h05130ba5_859307e0,
        64'h06130000_25170000,
        64'h2597b765_00979023,
        64'h43189381_8cf59301,
        64'h17821702_27910107,
        64'h871b16fd_6685405c,
        64'hf1718c2f_f0ef6585,
        64'h4681862e_84aebfc9,
        64'h0ee7ab23_47050000,
        64'h1797c03f_e0ef0f65,
        64'h051310a5_859307f0,
        64'h06130000_25170000,
        64'h25978082_610564a2,
        64'h644260e2_4505cb8d,
        64'h3037f793_439c9381,
        64'h17820247_879b415c,
        64'h02f71163_842a1117,
        64'h87931111_17b71407,
        64'ha2235158_00001797,
        64'hc541e426_e822ec06,
        64'h1101b6c1_4905ea05,
        64'h01e31f80_00ef8522,
        64'hb6f94905_eaf708e3,
        64'h47890b94_c703b5c1,
        64'hc4079de3_0a24c783,
        64'h00e78e63_4711bcd7,
        64'h13e30b94_c703bd39,
        64'h02f40e23_4785d85f,
        64'he0ef00e7_90230047,
        64'h67133e80_05130007,
        64'hd703b901_4905def7,
        64'h09e34785_0b94c703,
        64'hbe051ce3_285000ef,
        64'h852285a6_c00512e3,
        64'h688000ef_8522d47c,
        64'h4795bfd5_93411742,
        64'h0007d703_eb158b09,
        64'h93411742_0007d703,
        64'h00e79023_00176713,
        64'h0007d703_93811782,
        64'h02c7879b_c2070ee3,
        64'h8b210007_57039301,
        64'h170203e7_871b405c,
        64'hdfffe0ef_00e79023,
        64'h00876713_0007d703,
        64'h00e69023_93819341,
        64'h17429b69_93411742,
        64'h178203e7_879b0006,
        64'hd7039281_168202c7,
        64'h869b3885_05136505,
        64'h405cec07_9ee303c4,
        64'h4783eef7_12e347a1,
        64'h4858eee7_f6e3478d,
        64'h00d14703_bfbdd47c,
        64'h4795fee7_f5e34785,
        64'h03744703_dbed8b89,
        64'hbba1d3f1_0a24c783,
        64'hd47c4799_c71900c7,
        64'hf713b755_d47c4791,
        64'h00f9f863_03744783,
        64'hc30d00c7_f713b311,
        64'h892ab321_4905ee05,
        64'h05e34930_00ef8522,
        64'h10058593_03a205b7,
        64'hee079ee3_0a24c783,
        64'h12e6fb63_4685ffc7,
        64'h871b14e7_8c63471d,
        64'h547cd005_19e339f0,
        64'h00ef8522_85a6d005,
        64'h1fe37a20_00ef8522,
        64'hd47c479d_06e9f363,
        64'h03744703_cf210307,
        64'hf7130c44_c783d07c,
        64'h8fd90d44_c703d07c,
        64'h8fd90087_171b0d54,
        64'hc703d07c_27818fd9,
        64'h0107979b_0d64c783,
        64'hd0780187_971b0d74,
        64'hc783d605_15e33f70,
        64'h00ef1304_84938522,
        64'h13048593_00001497,
        64'hd80510e3_3da000ef,
        64'h8522bb45_4905d941,
        64'h011000ef_8522d47c,
        64'h4795f8e7_ffe34785,
        64'h03744703_d3dd8b89,
        64'h00d14783_d7dd0004,
        64'hc7831007_c9630024,
        64'h8783ed69_5ec000ef,
        64'h8522858a_dc0512e3,
        64'h41e000ef_8522c791,
        64'h8b910014_c783dc05,
        64'h1be33020_00ef8522,
        64'h85a6de05_11e33c30,
        64'h00ef8522_bd09e8f7,
        64'h08e34785_03444703,
        64'he8f71de3_47915478,
        64'h1efa6963_03744783,
        64'hc7898b89_0c44c783,
        64'hd07c8fd9_0d44c703,
        64'hd07c8fd9_0087171b,
        64'h0d54c703_d07c2781,
        64'h8fd90107_979b0d64,
        64'hc783d078_0187971b,
        64'h0d74c783_e2051ee3,
        64'h4c9000ef_20248493,
        64'h85222024_85930000,
        64'h1497e405_19e34ac0,
        64'h00ef8522_ef3a1be3,
        64'h03644a03_eee7ffe3,
        64'h478d0354_4703bdd9,
        64'hac058593_dc1c0121,
        64'hf5b7ac07_879b0121,
        64'hf7b7bf85_02f40a23,
        64'h4789bdcd_84058593,
        64'hdc1c017d_85b78407,
        64'h879b017d_87b702f7,
        64'h00634789_03644703,
        64'hea0514e3_de6ff0ef,
        64'h8522f0d7_11e3bdf1,
        64'h4905f0f7_05e34795,
        64'h00f6f763_0ff7f793,
        64'hfff7079b_46850344,
        64'h4703ffed_8b890007,
        64'h47839301_170202f7,
        64'h071b4058_00e78023,
        64'h47099381_00d71023,
        64'h17823ff6_869b9301,
        64'h76fd02f7_879b1702,
        64'h00c69023_0327871b,
        64'h92811682_0307869b,
        64'h567d405c_02f40a23,
        64'h4785c949_cb4ff0ef,
        64'h85221000_059340ff,
        64'h86374681_bf894905,
        64'h4ee7a723_47050000,
        64'h1797ffbf_e0ef4ee5,
        64'h05134ea5_859323f0,
        64'h06130000_25170000,
        64'h2597bfa5_00a03933,
        64'h3c2000ef_85222000,
        64'h0593f8f7_05e34791,
        64'h54781ee7_82634715,
        64'h10e78363_47091937,
        64'h87634985_03444783,
        64'hfd3d892a_d1cff0ef,
        64'h85227000_05934681,
        64'h4830f941_0e7000ef,
        64'h8522a805_8593dc1c,
        64'h018cc5b7_a807879b,
        64'h018cc7b7_f54dd55f,
        64'hf0ef8522_02f50a23,
        64'h4795fae7_91e38ff5,
        64'h40000737_c00006b7,
        64'h551c8082_610d7a46,
        64'h79e6690a_64aa854a,
        64'h644a60ea_490558e7,
        64'hae234705_00001797,
        64'h8a8ff0ef_59c50513,
        64'h59858593_24000613,
        64'h00002517_00002597,
        64'ha01d4905_cd69d9ef,
        64'hf0ef8522_45814601,
        64'h46819c0f_f0ef7105,
        64'h05136509_04f70b63,
        64'h47890205_0e23dd1c,
        64'ha807879b_000627b7,
        64'h03654703_02f50a23,
        64'h02f50ba3_478504f7,
        64'h1163842a_11178793,
        64'h111117b7_6007a523,
        64'h51580000_17971005,
        64'h0463fc02_f802f402,
        64'hf002ec02_e802e402,
        64'he0020004_b0239881,
        64'hf8d2fcce_e14ae922,
        64'hed0605f1_0493e526,
        64'h7135b5f1_d07c02e4,
        64'h0aa30097_d79b00f6,
        64'hf7130126_569b00e7,
        64'h97bb00f6_f71300e7,
        64'h97bb2785_0086d69b,
        64'h27098b1d_8fcd4210,
        64'h0077571b_8fe59201,
        64'h0167559b_160200a6,
        64'h979b2681_270101c7,
        64'h861b4294_43184210,
        64'h92819301_92011682,
        64'h17021602_0187869b,
        64'h0147871b_0107861b,
        64'hc0048493_405cf005,
        64'h15e3e8af_f0ef8522,
        64'h90048593_46816485,
        64'h4830fd11_e9cff0ef,
        64'h30000593_12340637,
        64'hc83cc438_123407b7,
        64'hc47cc070_c02c0007,
        64'hd7830007_57030006,
        64'h56030005_d5839381,
        64'h93019201_91811782,
        64'h17021602_158227f1,
        64'h0187871b_0147861b,
        64'h0107859b_85224681,
        64'h405cf535_eecff0ef,
        64'h85222000_05934601,
        64'h4681d81c_47850007,
        64'h54630217_97138082,
        64'h61054505_64a272e7,
        64'haa234705_00001797,
        64'h644260e2_a44ff0ef,
        64'h73850513_73458593,
        64'h67000613_00002517,
        64'h00002597_b751f6e7,
        64'h98e38ff5_40000737,
        64'hc00006b7_551c8082,
        64'h610564a2_644260e2,
        64'h450576e7_ac234705,
        64'h00001797_a84ff0ef,
        64'h77850513_77458593,
        64'h67100613_00002517,
        64'h00002597_80826105,
        64'h450564a2_644260e2,
        64'hd165f82f_f0ef8522,
        64'h10000593_40ff8637,
        64'h46810807_c8632781,
        64'h439c9381_178227c1,
        64'h405ca015_c911fa6f,
        64'hf0ef8522_45814601,
        64'h46810207_5b6302f7,
        64'h9713439c_93811782,
        64'h0247879b_405ccb99,
        64'h445c08f7_04634789,
        64'h03654703_06f71263,
        64'h842a1117_87931111,
        64'h17b78007_a4235158,
        64'h00002797_cd4de426,
        64'he822ec06_11018082,
        64'h61454501_69a26942,
        64'h64e200f6_90234789,
        64'h740270a2_b775dd25,
        64'h811ff0ef_84e79423,
        64'h85228005_8593864e,
        64'h4685470d_00002797,
        64'h6589b799_f4c713e3,
        64'h01077733_40000637,
        64'hc0000837_5518bff9,
        64'hf4064fe3_02f71613,
        64'h43189301_17020247,
        64'h871b8082_61454505,
        64'h69a26942_64e27402,
        64'h70a200f6_10233ff7,
        64'h879b9201_77fd1602,
        64'h0326061b_fe0756e3,
        64'h8b894107_571b0107,
        64'h971b93c1_17c20006,
        64'hd783e3c1_a0119281,
        64'h16820306_069b4050,
        64'hed0589bf_f0ef8ce7,
        64'h9a238522_90058593,
        64'h864e86a6_02700713,
        64'h00002797_658908f4,
        64'h88634785_dffff0ef,
        64'h852285a6_864ae13d,
        64'h79a000ef_20000593,
        64'h00f70763_842a89ae,
        64'h89362000_0713439c,
        64'h93811782_2791eb59,
        64'h45580ae8_0863415c,
        64'h84b24709_03654803,
        64'he44ee84a_f022f406,
        64'hec267179_80826145,
        64'h4501421c_69a26942,
        64'h64e29201_00f69023,
        64'h16024789_26417402,
        64'h70a2b775_dd25927f,
        64'hf0ef94e7_9f238522,
        64'h10058593_864e4685,
        64'h474d0000_27976585,
        64'hb799f4c7_13e30107,
        64'h77334000_0637c000,
        64'h08375518_bff9f406,
        64'h4fe302f7_16134318,
        64'h93011702_0247871b,
        64'h80826145_450569a2,
        64'h694264e2_740270a2,
        64'h00f61023_3ff7879b,
        64'h920177fd_16020326,
        64'h061bfe07_56e38b89,
        64'h4107571b_0107971b,
        64'h93c117c2_0006d783,
        64'he3c1a011_92811682,
        64'h0306069b_4050ed05,
        64'h9b1ff0ef_9ee79523,
        64'h85222005_8593864e,
        64'h86a60370_07130000,
        64'h27976585_08f48863,
        64'h4785f15f_f0ef8522,
        64'h85a6864a_e13d0b10,
        64'h00ef2000_059300f7,
        64'h0763842a_89ae8936,
        64'h20000713_439c9381,
        64'h17822791_eb594558,
        64'h0ae80863_415c84b2,
        64'h47090365_4803e44e,
        64'he84af022_f406ec26,
        64'h71798082_00a8a023,
        64'h08b79123_0208d893,
        64'h0805051b_08e79023,
        64'h08c7a223_18820230,
        64'h071397aa_0588889b,
        64'h83f50206_97930265,
        64'h85bb9e39_01e7073b,
        64'h7741ff07_18e307a1,
        64'h00ee073b_00079123,
        64'h01d79023_c3d86e41,
        64'h02100e93_873201e8,
        64'h083b0805_079300c8,
        64'h083b0107_1f1b7841,
        64'hce85fff7_069b0016,
        64'h871bc399_0006871b,
        64'h93c117c2_0107d69b,
        64'h04e86963_0007881b,
        64'h468102b3_07bb00f3,
        64'h73332601_67410007,
        64'hd7839381_17820048,
        64'h879b137d_63050045,
        64'h28838082_014100a0,
        64'h353360a2_acdff0ef,
        64'he4067000_05934681,
        64'h11414930_b339d07c,
        64'h0097d79b_00f717bb,
        64'h00f67793_00f7173b,
        64'h0086561b_27052789,
        64'h8b9d8f55_0077d79b,
        64'h8f650167_d69bc004,
        64'h849300a6_171bb381,
        64'hd07c00a7_979b2785,
        64'h93a9178a_d4d718e3,
        64'h4685cb19_8b0d0166,
        64'hd71b2601_0007079b,
        64'h43944290_43189301,
        64'h93819281_42101782,
        64'h16821702_920127f1,
        64'h16020187_869b0147,
        64'h871b0107_861b405c,
        64'hd4051be3_b5dff0ef,
        64'h85229004_85934681,
        64'h6485b599_02f40aa3,
        64'h4789bb85_4505d16d,
        64'hb79ff0ef_85223000,
        64'h05934601_4681ee19,
        64'hc8308e65_43909381,
        64'h178227c1_405ca809,
        64'hc47cc438_c074c030,
        64'h0007d783_00075703,
        64'h0006d683_00065603,
        64'h93819301_92819201,
        64'h17821702_16821602,
        64'h27f10187_871b0147,
        64'h869b0107_861b74c1,
        64'h405cdc05_18e3bd7f,
        64'hf0ef8522_20000593,
        64'h46014681_de0491e3,
        64'hfed79ee3_8ff1431c,
        64'h00d78663_8ff1431c,
        64'h93011702_0247071b,
        64'h01f006b7_01f00637,
        64'h4058821f_f0ef00f7,
        64'h10230047_e7933e80,
        64'h05130007_5783dfed,
        64'h8b890007_578300f7,
        64'h10230017_e7930007,
        64'h57839301_02079713,
        64'h02c7879b_e2070de3,
        64'h8b210007_57039301,
        64'h170203e7_871b405c,
        64'h867ff0ef_00f69023,
        64'h0087e793_38850513,
        64'h65050006_d7839281,
        64'h00f71023_93c117c2,
        64'h9be993c1_17c21682,
        64'h03e6869b_00075783,
        64'h93011702_02c6871b,
        64'hfff58ff1_431cc781,
        64'h8ff1431c_93011702,
        64'h0246871b_84aa01f0,
        64'h06374054_ca5ff0ef,
        64'h8522b005_85934601,
        64'h468102f4_0e236585,
        64'h47850c07_5d630277,
        64'h9713d818_47050007,
        64'h54630217_9713bf75,
        64'h41ff8637_fd4792e3,
        64'h485cfd37_95e340ff,
        64'h86378522_03644783,
        64'hee0513e3_85a64681,
        64'hcf1ff0ef_85224601,
        64'h85ca4681_0207c963,
        64'h2781439c_93811782,
        64'h27c1405c_f00515e3,
        64'hd11ff0ef_a8299004,
        64'h84934a21_49897009,
        64'h091364ad_690d02f4,
        64'h0aa34785_1af70f63,
        64'h1aa00713_431c9301,
        64'h17022741_40588082,
        64'h61454505_6a0269a2,
        64'h694264e2_d6e7a923,
        64'h47050000_27977402,
        64'h70a2883f_f0efd765,
        64'h0513d725_85931610,
        64'h06130000_35170000,
        64'h3597b785_f4e796e3,
        64'h8ff54000_0737c000,
        64'h06b7551c_a0a9ffed,
        64'h8b890006_c7839281,
        64'h168202f7_069b4058,
        64'h00a78023_93811782,
        64'h02f7879b_405cfaf5,
        64'h12e34789_c925daff,
        64'hf0ef8522_80058593,
        64'h1aa00613_46816585,
        64'h80826145_6a0269a2,
        64'h694264e2_740270a2,
        64'h4505dee7_ac234705,
        64'h00002797_905ff0ef,
        64'hdf850513_df458593,
        64'h16200613_00003517,
        64'h00003597_80826145,
        64'h6a0269a2_694264e2,
        64'h740270a2_4505c521,
        64'he09ff0ef_85224581,
        64'h46014681_00075963,
        64'h02f79713_439c9381,
        64'h17820247_879b405c,
        64'hcb99445c_0af70663,
        64'h4789c95c_47910365,
        64'h470304f7_1563842a,
        64'h11178793_111117b7,
        64'he607a723_51580000,
        64'h2797c16d_e052e44e,
        64'he84aec26_f022f406,
        64'h7179b769_00e79023,
        64'h25013ff7_071b777d,
        64'h4509e311_ffe57713,
        64'h91411542_0007d503,
        64'h93810205_17930325,
        64'h051b8082_61054505,
        64'h690264a2_eae7ad23,
        64'h47050000_27976442,
        64'h60e29cbf_f0efebe5,
        64'h0513eba5_859344b0,
        64'h06130000_35170000,
        64'h3597b76d_00f61023,
        64'h02000793_d6dd0206,
        64'hf6930006_56838082,
        64'h61056902_64a26442,
        64'h60e24505_f0e7a123,
        64'h47050000_2797a0ff,
        64'hf0eff025_0513efe5,
        64'h859344c0_06130000,
        64'h35170000_35978082,
        64'h61054501_690264a2,
        64'h00f61023_47856442,
        64'h60e2d7e5_0805c763,
        64'hc7318b85_4105d59b,
        64'h0107959b_93c117c2,
        64'h00065783_92011602,
        64'h0305061b_40c800a9,
        64'h20230209_59138d5d,
        64'h19028d75_29313fff,
        64'h06b70105_151bf767,
        64'hd7830000_2797efb5,
        64'h02057793_c7818b89,
        64'h439c9381_17820249,
        64'h079bcb19_25012701,
        64'hdff77713_9f21d007,
        64'h071b777d_e0bff0ef,
        64'h00e79023_93813ff7,
        64'h071b777d_178200d7,
        64'h10230329_079b9301,
        64'h17020309_071b0045,
        64'h2903c390_93811782,
        64'h27a1842e_56fd415c,
        64'h00e78023_47399381,
        64'h00d71023_17829301,
        64'h92c102e7_879b1702,
        64'h16c20067_871beb75,
        64'h8b054318_93011702,
        64'h0247871b_415c0ef7,
        64'h126384aa_11178793,
        64'h111117b7_0007a923,
        64'h51580000_27971405,
        64'h0063e04a_e426e822,
        64'hec061101_8082bdf9,
        64'h852ef4f5_85e3c007,
        64'h8793f8e5_8de31007,
        64'h8713f4f5_8de38082,
        64'h83a78513_eee68fe3,
        64'h81a78513_47050345,
        64'h46838082_31b00513,
        64'h808261b0_0513f0f7,
        64'h0ce363a0_05134785,
        64'h03454703_b715852e,
        64'hfcf58ce3_80078793,
        64'hf8d58ce3_40068693,
        64'hfee584e3_90078713,
        64'h6789feb7_71e3fee5,
        64'h8be37007_87138082,
        64'h03a5e513_f4f59ae3,
        64'h50078793_00e58663,
        64'h30078713_b78dfce5,
        64'h87e3d007_0713f6f5,
        64'h88e361a5_05136005,
        64'h07936521_8082f6f5,
        64'h9fe32090_05132000,
        64'h0793f8f5_86e31020,
        64'h05131000_07938082,
        64'h01a5e513_f8f59ee3,
        64'ha0078793_fae583e3,
        64'h90978513_90078713,
        64'h0ab76f63_00e58e63,
        64'hb0078713_8082fae5,
        64'h9fe39027_85139007,
        64'h8713fce5_86e333a7,
        64'h85133007_8713fce5,
        64'h8ce3a1a7_8513a007,
        64'h871367ad_06b7f663,
        64'h08f58c63_70070793,
        64'h67250ab7_746304e5,
        64'h8f637006_8713668d,
        64'h8082852e_12f58563,
        64'h51b00513_50000793,
        64'h00f58963_71a00513,
        64'h70000793_0ef58e63,
        64'h60000793_08b7f963,
        64'h10f58e63_30000793,
        64'h06b76c63_80078713,
        64'h12070963_8005871b,
        64'h04b76263_0ee58a63,
        64'h20078713_67858082,
        64'h01414505_1ae7a123,
        64'h47050000_27976402,
        64'h60a2cb3f_f0ef1a65,
        64'h05131a25_85930b50,
        64'h06130000_35170000,
        64'h35978082_01414505,
        64'h1ce7a723_47050000,
        64'h27976402_60a2cdff,
        64'hf0ef1d25_05131ce5,
        64'h85930b40_06130000,
        64'h35170000_3597b791,
        64'h472df406_d5e34705,
        64'h02579693_f406cae3,
        64'h47350267_9693b781,
        64'hdffff0ef_0c800513,
        64'hf4e796e3_8ff54000,
        64'h0737c000_06b7541c,
        64'h80820141_45056402,
        64'h60a2b709_00f60023,
        64'h47c18082_014100e7,
        64'h90232000_07139381,
        64'h24d71523_17820000,
        64'h271746cd_00071023,
        64'h27919301_00069023,
        64'h17029281_03a7871b,
        64'h168200c7_10233ff6,
        64'h061b0387_869b9301,
        64'h767d1702_00c69023,
        64'h0367871b_92811682,
        64'h0347869b_640260a2,
        64'h405c00e7_80239381,
        64'h17820287_879b4741,
        64'h405c00e7_80239381,
        64'h17820297_879beff0,
        64'h0613405c_0a06d563,
        64'h02779693_473d541c,
        64'he9416540_10ef8522,
        64'ha8058593_000625b7,
        64'h0af70663_47890364,
        64'h470300f6_80239281,
        64'hd41047bd_16820296,
        64'h869b4310_930102f4,
        64'h0b230ff7_f7931702,
        64'h0406871b_0007d783,
        64'h93811782_0fe6879b,
        64'hffed8b85_00074783,
        64'h93011702_02f6871b,
        64'h405400e7_80239381,
        64'h178202f7_879b4705,
        64'h405cf19f_f0ef3e80,
        64'h05130006_002310e7,
        64'h80639201_47090ff7,
        64'hf7930604_38230604,
        64'h22231602_d4780296,
        64'h061b4719_0007d783,
        64'h938102e4_00231782,
        64'h0fe6079b_0205c703,
        64'hcc58cc14_c8480104,
        64'h28230114_2623d05c,
        64'hc0500064_10231117,
        64'h879b1111_17b7c41c,
        64'h4d9449c8_0105a803,
        64'h00c5a883_0005d303,
        64'h4dd8842a_459c1c05,
        64'h8c633807_af230000,
        64'h27971a05_0c63e022,
        64'he4061141_8082f2e5,
        64'h05130000_25178082,
        64'hf5c50513_00002517,
        64'h808200e7_83634501,
        64'h0247d783_f4c78793,
        64'h00002797_02a78163,
        64'h872af5a7_d7830000,
        64'h27978082_fea7ede3,
        64'h8f99ff86_b7830200,
        64'hc6b702f5_05330280,
        64'h0793fee7_8ee3ff86,
        64'hb7030200_c6b7ff87,
        64'hb7830200_c7b78082,
        64'hff87b503_0200c7b7,
        64'h80826125_70a2a1bf,
        64'hf0efe43a_ecc6e8c2,
        64'he4bef406_72c50513,
        64'h567d080c_86b21838,
        64'hec2ee0ba_fc36ffff,
        64'hf517e82a_711da43f,
        64'hf06f72e5_0513ffff,
        64'hf51785aa_862e86b2,
        64'h87368082_610560e2,
        64'ha5dff0ef_ec06a645,
        64'h0513002c_567d872e,
        64'h00000517_86aa1101,
        64'h80826161_60e2a7bf,
        64'hf0efe43a_e4c6e0c2,
        64'hfc3eec06_10387745,
        64'h0513f83a_fffff517,
        64'h85aa862e_86b2f436,
        64'h715d8082_616160e2,
        64'haa5ff0ef_e43ae4c6,
        64'he0c2fc3e_ec067a25,
        64'h05131018_567df83a,
        64'hf032ffff_f51785aa,
        64'h86aef436_715d8082,
        64'h612560e2_ad1ff0ef,
        64'he43aecc6_e8c2e4be,
        64'hec06ae65_0513567d,
        64'h1038858a_e0baf832,
        64'hf42e0000_051786aa,
        64'hfc36711d_b31d4809,
        64'hb32d4821_bb1d4841,
        64'h0206e693_bb498da2,
        64'h99020250_051385d2,
        64'h866e86ce_001d8413,
        64'hb7d58622_2c859902,
        64'h00160413_02000513,
        64'h85d286ce_bb6d8db2,
        64'h8aea018c_e563c019,
        64'hfc089de3_fff8869b,
        64'hfe0a82e3_c51901b7,
        64'h06330007_450378a2,
        64'h77029902_85d286ce,
        64'hf83af03a_f4460705,
        64'h88b6b7e1_78c28df2,
        64'h8cc27762_7e027822,
        64'h99020200_051385d2,
        64'h86ce866e_f072f442,
        64'hf846fc3a_001d8e13,
        64'hb7c90785_a08140ed,
        64'h8db38cc2_018ce863,
        64'h001c881b_e4110006,
        64'h841b8a89_00060c9b,
        64'h8666011c_f3638646,
        64'h000a8863_40e78cbb,
        64'h2a814006_fa9302f6,
        64'h1b63c199_0007c583,
        64'h87ba00f7_06339381,
        64'h02089793_00088563,
        64'h57fd000a_b703008a,
        64'h8d13b7cd_8ca22b05,
        64'h99020200_051385d2,
        64'h86ce001c_84138666,
        64'hb5598de6_8aea018b,
        64'h6563c019_9902001d,
        64'h8c93008a_8d1385d2,
        64'h866e86ce_000ac503,
        64'hff8764e3_001d8d13,
        64'h00170b1b_8dea875a,
        64'h99020200_051385d2,
        64'h86ce866e_a8094705,
        64'he00d4b05_0006841b,
        64'h8a89b7ed_8f7d67e2,
        64'hdbe50807_f793b769,
        64'h93014781_e062e436,
        64'h17020ff7_7713ca09,
        64'h000aa703_0407f613,
        64'hb755e062_e4364781,
        64'h000ab703_c7191007,
        64'hf713bde5_4781e062,
        64'he436000a_b703c719,
        64'hbff1000a_a783b7cd,
        64'h000a9783_c7810807,
        64'hf793bfd9_40e6073b,
        64'h93fde062_e43600e7,
        64'hc63341f7_d71b000a,
        64'hc783cf09_0406f713,
        64'hb789bb7f_f0ef854a,
        64'h85d2866e_86ce93fd,
        64'h40e60733_00f74633,
        64'h43f7d713_e062e436,
        64'h000ab783_c31d87b6,
        64'h1006f713_b5dd0780,
        64'h0793eef5_09e30750,
        64'h0793a89d_4841e03e,
        64'he436008a_8413000a,
        64'hb70347c1_0216e693,
        64'hd4f51ae3_07000793,
        64'hf0f50ce3_06f00793,
        64'h02a7e563_12f50f63,
        64'h07300793_b71d0640,
        64'h07930ef5_06630630,
        64'h0793bddd_0c06e693,
        64'h8082614d_6da66d46,
        64'h6ce67c06_7ba67b46,
        64'h7ae66a0a_69aa694a,
        64'h64ea000d_851b740a,
        64'h70aa9902_450185d2,
        64'h86cefff9_8613013d,
        64'he463866e_da0517e3,
        64'h0004c503_8aa28daa,
        64'hcf5ff0ef_854a85d2,
        64'h866e86ce_93fd40e6,
        64'h073300f7_463343f7,
        64'hd713e062_e436000a,
        64'hb783cf45_10c51c63,
        64'h06400613_00c50663,
        64'h008a8413_02085813,
        64'h270187b6_06900613,
        64'h18022006_f7139af9,
        64'hc3914006_f7939acd,
        64'h00f50363_06400793,
        64'h00f50763_48299abd,
        64'h06900793_2ef50463,
        64'h06200793_2ef50663,
        64'h06f00793_2ef50663,
        64'h05800793_2ef50c63,
        64'h07800793_e4f514e3,
        64'h05800793_2ef50863,
        64'h02500793_0ca7ef63,
        64'h00f50c63_06200793,
        64'h0ea7ec63_02f50263,
        64'h00170493_06900793,
        64'h00074503_0806e693,
        64'h0ef60e63_0014c603,
        64'ha0390024_87133006,
        64'he693a821_1006e693,
        64'h00f60563_0014c603,
        64'hb7e907a0_061300c7,
        64'h89630740_0613bf65,
        64'h84babf75_8abe0489,
        64'h28814881_0008d363,
        64'h008a8793_000aa883,
        64'h00f61d63_02a00793,
        64'ha8998726_04c78063,
        64'h06a00613_04c78c63,
        64'h06800613_02f66d63,
        64'h04c78663_00148713,
        64'h06c00613_0004c783,
        64'hfef671e3_0ff7f793,
        64'hfd07079b_00148593,
        64'h0004c703_00e888bb,
        64'hfd08889b_84ae031b,
        64'h88bbb775_84b28aba,
        64'h40f00c3b_0026e693,
        64'h0007d663_00078c1b,
        64'h008a8713_000aa783,
        64'hfce796e3_4c0102a0,
        64'h0713a825_462584ba,
        64'h06f5ee63_4006e693,
        64'h0ff7f793_fd06079b,
        64'h00148713_45a50014,
        64'hc60306f7_17634881,
        64'h02e00793_0004c703,
        64'hfef671e3_0ff7f793,
        64'hfd07079b_00148593,
        64'h0004c703_00e30c3b,
        64'hfd03031b_84ae038b,
        64'h833bbf75_0106e693,
        64'hb7c90086_e693b7e1,
        64'h0046e693_b7f90026,
        64'he693a025_46254c01,
        64'h06e5e963_45a50ff7,
        64'h7713fd07_871b02a7,
        64'h856302b7_8463fcf7,
        64'h6fe302e7_85630014,
        64'h86130004_c78384b2,
        64'h0016e693_02879163,
        64'h03000413_02878f63,
        64'h02d00413_a8210230,
        64'h05130200_059302b0,
        64'h07134681_a15585d2,
        64'h866e86ce_001d8413,
        64'h00f50863_04850250,
        64'h0793ac81_4ba9ec3e,
        64'h4d81fffb_07936b41,
        64'hcc890913_00000917,
        64'he589892a_8aba84b6,
        64'h89b28a2e_e4eee8ea,
        64'hece6f0e2_f4def8da,
        64'hf122f506_fcd6e152,
        64'he54ee94a_ed267171,
        64'h80829a1f_f06fc119,
        64'hb7e1006e_033b8082,
        64'h616160a6_d17ff0ef,
        64'h887e1018_0008089b,
        64'he43ae876_e0464746,
        64'hfc579de3_c319fe6f,
        64'h0fa39f3e_0ff37313,
        64'h02010f13_07850307,
        64'h57330303_031b03e3,
        64'hee630fff_73130307,
        64'h7f330200_0293ff63,
        64'h0e1b43a5_47810410,
        64'h0313000e_04630610,
        64'h0313020e_fe13c721,
        64'h47810003_0463400e,
        64'hf313fefe_fe93e319,
        64'h4ee68fbe_e486715d,
        64'hb7e1006e_033b8082,
        64'h616160a6_d97ff0ef,
        64'h887e1018_0008089b,
        64'he43ae876_e0464746,
        64'hfc579de3_c319fe6f,
        64'h0fa39f3e_0ff37313,
        64'h02010f13_07850307,
        64'h57330303_031b03e3,
        64'hee630fff_73130307,
        64'h7f330200_0293ff63,
        64'h0e1b43a5_47810410,
        64'h0313000e_04630610,
        64'h0313020e_fe13c721,
        64'h47810003_0463400e,
        64'hf313fefe_fe93e319,
        64'h4ee68fbe_e486715d,
        64'hb7a98622_9b020016,
        64'h04130200_051385de,
        64'h86e2b791_9b0285de,
        64'h86e20009_4503b7ed,
        64'h41540cb3_02095913,
        64'h02099913_bf89ff27,
        64'he3e3009c_87b384ea,
        64'h00148d13_67229b02,
        64'he43a0200_051385de,
        64'h86e28626_b7ad00d6,
        64'h00230087_0633da3d,
        64'h0087f613_bf9d02b0,
        64'h06130087_06b3c611,
        64'h0047f613_bfa10620,
        64'h06130087_06b3f886,
        64'hece346fd_f6d898e3,
        64'h4689b7bd_05800613,
        64'h008706b3_fa86e7e3,
        64'h46fd8082_61658532,
        64'h6d426ce2_7c027ba2,
        64'h7b427ae2_6a0669a6,
        64'h694664e6_740670a6,
        64'h0b37e163_415607b3,
        64'h0209d993_1982000a,
        64'h09630094_06330b2c,
        64'h9663197d_412d0633,
        64'h01248d33_fff70c93,
        64'h00870933_cbcd84d6,
        64'h8b8d0405_00c68023,
        64'h02d00613_008706b3,
        64'h08080463_00d40b63,
        64'h02000693_040500c6,
        64'h80230300_06130087,
        64'h06b30286_e66346fd,
        64'h040500c6_80230780,
        64'h06130087_06b30486,
        64'he06346fd_ead10207,
        64'hf6930ad8_966346c1,
        64'h4401bf55_fe6e0fa3,
        64'h00870e33_0405a0e9,
        64'h02c89a63_84364609,
        64'h02c88163_14794641,
        64'hc285fff4_06930286,
        64'h95639281_02099693,
        64'h00868763_92811682,
        64'hcc0dee15_4007f613,
        64'hca3d0107_f61302b4,
        64'h1e6300a4_7463c609,
        64'h03000313_02000593,
        64'h91010209_9513fea4,
        64'h69e3fe6e_0fa30087,
        64'h0e330405_00b40963,
        64'ha8010300_03130200,
        64'h05939101_02069513,
        64'h39fdc191_00c7f593,
        64'h00081563_c6190009,
        64'h89630017_f613040a,
        64'h1a6359e6_56c68ab2,
        64'h8bae8b2a_8c362a01,
        64'he86aec66_e8caeca6,
        64'hf486f062_f45ef85a,
        64'hfc560027_fa13e4ce,
        64'he0d2478a_843ef0a2,
        64'h71598082_8302658c,
        64'h0005b303_c5098082,
        64'h808200a5_802395b2,
        64'h00d67563_bbe102f0,
        64'h00efd0a5_05130000,
        64'h4517bd35_ace50513,
        64'h85a60000_45170470,
        64'h00efac25_05130000,
        64'h4517cd09_84aadabf,
        64'hf0ef8552_865a020a,
        64'ha5830630_00efd265,
        64'h05130000_4517f579,
        64'h90e30804_84930770,
        64'h00ef2985_aac50513,
        64'h00004517_ff2c17e3,
        64'h089000ef_0905cc65,
        64'h05130000_45170009,
        64'h45830704_8c130284,
        64'h89130a30_00efd4e5,
        64'h05130000_45170af0,
        64'h00efd425_05130000,
        64'h4517708c_0bd000ef,
        64'hd3850513_00004517,
        64'h6c8c0cb0_00efd2e5,
        64'h05130000_4517688c,
        64'hff2c17e3_0dd000ef,
        64'h0905d1a5_05130000,
        64'h45170009_45830109,
        64'h0c130f30_00efd365,
        64'h05130000_4517fe99,
        64'h17e31030_00ef0905,
        64'hd4050513_00004517,
        64'h00094583_ff048913,
        64'h119000ef_d3450513,
        64'h00004517_125000ef,
        64'hd2a50513_85ce0000,
        64'h4517bf15_d1650513,
        64'h85ce0000_451713f0,
        64'h00efbba5_05130000,
        64'h4517cd09_4b910804,
        64'h89aa8a8a_ea9ff0ef,
        64'h850a4605_710144ac,
        64'h161000ef_d2450513,
        64'h00004517_45d616f0,
        64'h00efd125_05130000,
        64'h451745c6_17d000ef,
        64'hcf850513_00004517,
        64'h65a618b0_00efcee5,
        64'h05130000_45177582,
        64'h199000ef_ce450513,
        64'h00004517_65e21a70,
        64'h00efcda5_05130000,
        64'h451745d2_1b5000ef,
        64'hcd050513_00004517,
        64'h45c21c30_00efcc65,
        64'h05130000_451745b2,
        64'h1d1000ef_cbc50513,
        64'h00004517_45a21df0,
        64'h00efcb25_05130000,
        64'h45176582_1ed000ef,
        64'hca050513_00004517,
        64'hb75554f9_1fd000ef,
        64'hc9050513_00004517,
        64'hfa843583_20d000ef,
        64'hc8850513_00004517,
        64'hfaa43423_c11df73f,
        64'hf0ef848a_850a4585,
        64'h46057101_22d000ef,
        64'hc9050513_00004517,
        64'h80826125_6c426be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_64468526,
        64'h60e6fa04_011354fd,
        64'h259000ef_c9450513,
        64'h00004517_c51df4df,
        64'hf0ef8b2e_8a2a1080,
        64'he862ec5e_f456fc4e,
        64'he0cae4a6_ec86f05a,
        64'hf852e8a2_711d8082,
        64'h014160a2_557d28f0,
        64'h00efcb25_05130000,
        64'h4517c901_55e010ef,
        64'he406c1e5_05134605,
        64'h11410000_351786aa,
        64'hbfc94501_2b5000ef,
        64'hcb850513_00004517,
        64'hb7cd5575_2c5000ef,
        64'hca850513_00004517,
        64'hc90914c0_10ef8522,
        64'h80820141_640260a2,
        64'h55792e30_00efcae5,
        64'h05130000_4517cd01,
        64'h441000ef_8522c704,
        64'h041341d0_00003417,
        64'hc18d557d_85aa4210,
        64'h00ef4501_30d000ef,
        64'he022e406_cc650513,
        64'h11410000_45178082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_00a78223,
        64'h0ff57513_00d78023,
        64'h0085551b_0ff57693,
        64'h00d78623_f8000693,
        64'h00078223_01e71793,
        64'h470d02b5_553b0045,
        64'h959b8082_00a78023,
        64'hdf650207_77130147,
        64'hc70307fa_478d8082,
        64'h02057513_0147c503,
        64'h07fa478d_80820005,
        64'h45038082_00b50023,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_100004b7,
        64'h18858593_00003597,
        64'hf1402573_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_3d3020ef,
        64'h40000137_03249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
