/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 1151;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd0080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h08090000_38000000,
        64'hda0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha0018402_14458593,
        64'h00000597_10000437,
        64'he901c16f_f0ef1000,
        64'h053765a1_effff0ef,
        64'hd4050513_00001517,
        64'hd95fe0ef_e406a005,
        64'h05132005_85931141,
        64'h02626537_65f18082,
        64'h612570a2_a1bff0ef,
        64'he43aecc6_e8c2e4be,
        64'hf40672c5_0513567d,
        64'h080c86b2_1838ec2e,
        64'he0bafc36_fffff517,
        64'he82a711d_a43ff06f,
        64'h72e50513_fffff517,
        64'h85aa862e_86b28736,
        64'h80826105_60e2a5df,
        64'hf0efec06_a6450513,
        64'h002c567d_872e0000,
        64'h051786aa_11018082,
        64'h616160e2_a7bff0ef,
        64'he43ae4c6_e0c2fc3e,
        64'hec061038_77450513,
        64'hf83affff_f51785aa,
        64'h862e86b2_f436715d,
        64'h80826161_60e2aa5f,
        64'hf0efe43a_e4c6e0c2,
        64'hfc3eec06_7a250513,
        64'h1018567d_f83af032,
        64'hfffff517_85aa86ae,
        64'hf436715d_80826125,
        64'h60e2ad1f_f0efe43a,
        64'hecc6e8c2_e4beec06,
        64'hae650513_567d1038,
        64'h858ae0ba_f832f42e,
        64'h00000517_86aafc36,
        64'h711db31d_4809b32d,
        64'h4821bb1d_48410206,
        64'he693bb49_8da29902,
        64'h02500513_85d2866e,
        64'h86ce001d_8413b7d5,
        64'h86222c85_99020016,
        64'h04130200_051385d2,
        64'h86cebb6d_8db28aea,
        64'h018ce563_c019fc08,
        64'h9de3fff8_869bfe0a,
        64'h82e3c519_01b70633,
        64'h00074503_78a27702,
        64'h990285d2_86cef83a,
        64'hf03af446_070588b6,
        64'hb7e178c2_8df28cc2,
        64'h77627e02_78229902,
        64'h02000513_85d286ce,
        64'h866ef072_f442f846,
        64'hfc3a001d_8e13b7c9,
        64'h0785a081_40ed8db3,
        64'h8cc2018c_e863001c,
        64'h881be411_0006841b,
        64'h8a890006_0c9b8666,
        64'h011cf363_8646000a,
        64'h886340e7_8cbb2a81,
        64'h4006fa93_02f61b63,
        64'hc1990007_c58387ba,
        64'h00f70633_93810208,
        64'h97930008_856357fd,
        64'h000ab703_008a8d13,
        64'hb7cd8ca2_2b059902,
        64'h02000513_85d286ce,
        64'h001c8413_8666b559,
        64'h8de68aea_018b6563,
        64'hc0199902_001d8c93,
        64'h008a8d13_85d2866e,
        64'h86ce000a_c503ff87,
        64'h64e3001d_8d130017,
        64'h0b1b8dea_875a9902,
        64'h02000513_85d286ce,
        64'h866ea809_4705e00d,
        64'h4b050006_841b8a89,
        64'hb7ed8f7d_67e2dbe5,
        64'h0807f793_b7699301,
        64'h4781e062_e4361702,
        64'h0ff77713_ca09000a,
        64'ha7030407_f613b755,
        64'he062e436_4781000a,
        64'hb703c719_1007f713,
        64'hbde54781_e062e436,
        64'h000ab703_c719bff1,
        64'h000aa783_b7cd000a,
        64'h9783c781_0807f793,
        64'hbfd940e6_073b93fd,
        64'he062e436_00e7c633,
        64'h41f7d71b_000ac783,
        64'hcf090406_f713b789,
        64'hbb7ff0ef_854a85d2,
        64'h866e86ce_93fd40e6,
        64'h073300f7_463343f7,
        64'hd713e062_e436000a,
        64'hb783c31d_87b61006,
        64'hf713b5dd_07800793,
        64'heef509e3_07500793,
        64'ha89d4841_e03ee436,
        64'h008a8413_000ab703,
        64'h47c10216_e693d4f5,
        64'h1ae30700_0793f0f5,
        64'h0ce306f0_079302a7,
        64'he56312f5_0f630730,
        64'h0793b71d_06400793,
        64'h0ef50663_06300793,
        64'hbddd0c06_e6938082,
        64'h614d6da6_6d466ce6,
        64'h7c067ba6_7b467ae6,
        64'h6a0a69aa_694a64ea,
        64'h000d851b_740a70aa,
        64'h99024501_85d286ce,
        64'hfff98613_013de463,
        64'h866eda05_17e30004,
        64'hc5038aa2_8daacf5f,
        64'hf0ef854a_85d2866e,
        64'h86ce93fd_40e60733,
        64'h00f74633_43f7d713,
        64'he062e436_000ab783,
        64'hcf4510c5_1c630640,
        64'h061300c5_0663008a,
        64'h84130208_58132701,
        64'h87b60690_06131802,
        64'h2006f713_9af9c391,
        64'h4006f793_9acd00f5,
        64'h03630640_079300f5,
        64'h07634829_9abd0690,
        64'h07932ef5_04630620,
        64'h07932ef5_066306f0,
        64'h07932ef5_06630580,
        64'h07932ef5_0c630780,
        64'h0793e4f5_14e30580,
        64'h07932ef5_08630250,
        64'h07930ca7_ef6300f5,
        64'h0c630620_07930ea7,
        64'hec6302f5_02630017,
        64'h04930690_07930007,
        64'h45030806_e6930ef6,
        64'h0e630014_c603a039,
        64'h00248713_3006e693,
        64'ha8211006_e69300f6,
        64'h05630014_c603b7e9,
        64'h07a00613_00c78963,
        64'h07400613_bf6584ba,
        64'hbf758abe_04892881,
        64'h48810008_d363008a,
        64'h8793000a_a88300f6,
        64'h1d6302a0_0793a899,
        64'h872604c7_806306a0,
        64'h061304c7_8c630680,
        64'h061302f6_6d6304c7,
        64'h86630014_871306c0,
        64'h06130004_c783fef6,
        64'h71e30ff7_f793fd07,
        64'h079b0014_85930004,
        64'hc70300e8_88bbfd08,
        64'h889b84ae_031b88bb,
        64'hb77584b2_8aba40f0,
        64'h0c3b0026_e6930007,
        64'hd6630007_8c1b008a,
        64'h8713000a_a783fce7,
        64'h96e34c01_02a00713,
        64'ha8254625_84ba06f5,
        64'hee634006_e6930ff7,
        64'hf793fd06_079b0014,
        64'h871345a5_0014c603,
        64'h06f71763_488102e0,
        64'h07930004_c703fef6,
        64'h71e30ff7_f793fd07,
        64'h079b0014_85930004,
        64'hc70300e3_0c3bfd03,
        64'h031b84ae_038b833b,
        64'hbf750106_e693b7c9,
        64'h0086e693_b7e10046,
        64'he693b7f9_0026e693,
        64'ha0254625_4c0106e5,
        64'he96345a5_0ff77713,
        64'hfd07871b_02a78563,
        64'h02b78463_fcf76fe3,
        64'h02e78563_00148613,
        64'h0004c783_84b20016,
        64'he6930287_91630300,
        64'h04130287_8f6302d0,
        64'h0413a821_02300513,
        64'h02000593_02b00713,
        64'h4681a155_85d2866e,
        64'h86ce001d_841300f5,
        64'h08630485_02500793,
        64'hac814ba9_ec3e4d81,
        64'hfffb0793_6b41cc89,
        64'h09130000_0917e589,
        64'h892a8aba_84b689b2,
        64'h8a2ee4ee_e8eaece6,
        64'hf0e2f4de_f8daf122,
        64'hf506fcd6_e152e54e,
        64'he94aed26_71718082,
        64'hcc4ff06f_c119b7e1,
        64'h006e033b_80826161,
        64'h60a6d17f_f0ef887e,
        64'h10180008_089be43a,
        64'he876e046_4746fc57,
        64'h9de3c319_fe6f0fa3,
        64'h9f3e0ff3_73130201,
        64'h0f130785_03075733,
        64'h0303031b_03e3ee63,
        64'h0fff7313_03077f33,
        64'h02000293_ff630e1b,
        64'h43a54781_04100313,
        64'h000e0463_06100313,
        64'h020efe13_c7214781,
        64'h00030463_400ef313,
        64'hfefefe93_e3194ee6,
        64'h8fbee486_715db7e1,
        64'h006e033b_80826161,
        64'h60a6d97f_f0ef887e,
        64'h10180008_089be43a,
        64'he876e046_4746fc57,
        64'h9de3c319_fe6f0fa3,
        64'h9f3e0ff3_73130201,
        64'h0f130785_03075733,
        64'h0303031b_03e3ee63,
        64'h0fff7313_03077f33,
        64'h02000293_ff630e1b,
        64'h43a54781_04100313,
        64'h000e0463_06100313,
        64'h020efe13_c7214781,
        64'h00030463_400ef313,
        64'hfefefe93_e3194ee6,
        64'h8fbee486_715db7a9,
        64'h86229b02_00160413,
        64'h02000513_85de86e2,
        64'hb7919b02_85de86e2,
        64'h00094503_b7ed4154,
        64'h0cb30209_59130209,
        64'h9913bf89_ff27e3e3,
        64'h009c87b3_84ea0014,
        64'h8d136722_9b02e43a,
        64'h02000513_85de86e2,
        64'h8626b7ad_00d60023,
        64'h00870633_da3d0087,
        64'hf613bf9d_02b00613,
        64'h008706b3_c6110047,
        64'hf613bfa1_06200613,
        64'h008706b3_f886ece3,
        64'h46fdf6d8_98e34689,
        64'hb7bd0580_06130087,
        64'h06b3fa86_e7e346fd,
        64'h80826165_85326d42,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a60b37,
        64'he1634156_07b30209,
        64'hd9931982_000a0963,
        64'h00940633_0b2c9663,
        64'h197d412d_06330124,
        64'h8d33fff7_0c930087,
        64'h0933cbcd_84d68b8d,
        64'h040500c6_802302d0,
        64'h06130087_06b30808,
        64'h046300d4_0b630200,
        64'h06930405_00c68023,
        64'h03000613_008706b3,
        64'h0286e663_46fd0405,
        64'h00c68023_07800613,
        64'h008706b3_0486e063,
        64'h46fdead1_0207f693,
        64'h0ad89663_46c14401,
        64'hbf55fe6e_0fa30087,
        64'h0e330405_a0e902c8,
        64'h9a638436_460902c8,
        64'h81631479_4641c285,
        64'hfff40693_02869563,
        64'h92810209_96930086,
        64'h87639281_1682cc0d,
        64'hee154007_f613ca3d,
        64'h0107f613_02b41e63,
        64'h00a47463_c6090300,
        64'h03130200_05939101,
        64'h02099513_fea469e3,
        64'hfe6e0fa3_00870e33,
        64'h040500b4_0963a801,
        64'h03000313_02000593,
        64'h91010206_951339fd,
        64'hc19100c7_f5930008,
        64'h1563c619_00098963,
        64'h0017f613_040a1a63,
        64'h59e656c6_8ab28bae,
        64'h8b2a8c36_2a01e86a,
        64'hec66e8ca_eca6f486,
        64'hf062f45e_f85afc56,
        64'h0027fa13_e4cee0d2,
        64'h478a843e_f0a27159,
        64'h80828302_658c0005,
        64'hb303c509_80828082,
        64'h00a58023_95b200d6,
        64'h7563bbb5_efcff0ef,
        64'h97850513_00002517,
        64'hb3f56d25_05130000,
        64'h1517f94f_f0ef8526,
        64'hf18ff0ef_7d450513,
        64'h00001517_f24ff0ef,
        64'h7c850513_00001517,
        64'hc50d84aa_c33ff0ef,
        64'h8552865a_020aa583,
        64'hf40ff0ef_9a450513,
        64'h00002517_f57993e3,
        64'h08048493_f54ff0ef,
        64'h29857225_05130000,
        64'h1517ff2c_1be382bf,
        64'hf0ef0905_00094503,
        64'hf70ff0ef_9c450513,
        64'h00002517_ffeff0ef,
        64'h7088f82f_f0ef9c65,
        64'h05130000_2517811f,
        64'hf0ef6c88_f94ff0ef,
        64'h9c850513_00002517,
        64'h823ff0ef_07048c13,
        64'h02848913_6888faef,
        64'hf0ef9d25_05130000,
        64'h2517ff2c_1be3883f,
        64'hf0ef0905_00094503,
        64'h01090c13_fccff0ef,
        64'h9d050513_00002517,
        64'hfe991be3_8a1ff0ef,
        64'h09050009_4503ff04,
        64'h8913feaf_f0ef9ce5,
        64'h05130000_25178bbf,
        64'hf0ef0ff9_f513ffef,
        64'hf0ef9ca5_05130000,
        64'h2517b5fd_7d450513,
        64'h00001517_897ff0ef,
        64'h854e81bf_f0ef8d65,
        64'h05130000_2517827f,
        64'hf0ef8ca5_05130000,
        64'h2517c50d_080489aa,
        64'h8a8ad39f_f0ef850a,
        64'h46057101_04892583,
        64'h849ff0ef_81450513,
        64'h00002517_897ff0ef,
        64'h455685bf_f0efa065,
        64'h05130000_25178a9f,
        64'hf0ef4546_86dff0ef,
        64'h9f850513_00002517,
        64'h8fbff0ef_652687ff,
        64'hf0ef9ea5_05130000,
        64'h251790df_f0ef7502,
        64'h891ff0ef_9ec50513,
        64'h00002517_91fff0ef,
        64'h65628a3f_f0ef9e65,
        64'h05130000_25178f1f,
        64'hf0ef4552_8b5ff0ef,
        64'h9e850513_00002517,
        64'h903ff0ef_45428c7f,
        64'hf0ef9ea5_05130000,
        64'h2517915f_f0ef4532,
        64'h8d9ff0ef_9ec50513,
        64'h00002517_927ff0ef,
        64'h45228ebf_f0ef9ee5,
        64'h05130000_2517979f,
        64'hf0ef4b91_65028fff,
        64'hf0ef9f25_05130000,
        64'h251790bf_f0ef9de5,
        64'h05130000_2517bf61,
        64'h54f991bf_f0ef8e65,
        64'h05130000_25179a9f,
        64'hf0ef8526_92dff0ef,
        64'h9e850513_00002517,
        64'h939ff0ef_9dc50513,
        64'h00002517_c90584aa,
        64'h890ae49f_f0ef850a,
        64'h45854605_7101957f,
        64'hf0ef9e25_05130000,
        64'h25178082_61616c02,
        64'h6ba26b42_6ae27a02,
        64'h79a27942_74e26406,
        64'h852660a6_fb040113,
        64'h54fd983f_f0ef9e65,
        64'h05130000_2517c51d,
        64'hdf3ff0ef_8b2e8a2a,
        64'h0880e062_e45eec56,
        64'hf44ef84a_fc26e486,
        64'he85af052_e0a2715d,
        64'hb7655479_80826169,
        64'h6baa6b4a_6aea7a0a,
        64'h79aa794a_74ea640e,
        64'h60ae8522_547d9cff,
        64'hf0efa0a5_05130000,
        64'h2517c59f_f0efc5df,
        64'hf0efc61f_f0efc65f,
        64'hf0efc69f_f0efc6df,
        64'hf0efc71f_f0efc75f,
        64'hf0efa805_c7bff0ef,
        64'hc87ff0ef_45314581,
        64'h46054401_f93046e3,
        64'h19fda13f_f0efa6e5,
        64'h05130000_2517e799,
        64'h0359e7b3_07241a63,
        64'h29019041_14428c49,
        64'hcafff0ef_90410305,
        64'h141384a2_0085151b,
        64'hcbfff0ef_fd641ae3,
        64'h04040413_ff7497e3,
        64'h892af13f_f0ef0485,
        64'h854a0007_c5830094,
        64'h07b30400_0b934481,
        64'hc67ff0ef_850a0400,
        64'h05938622_49018426,
        64'h20048b13_ff451ee3,
        64'hcffff0ef_3e800a93,
        64'h0fe00a13_e951d15f,
        64'hf0ef4549_85a20ff6,
        64'h76130016_66130015,
        64'h161bf49f_f0ef0ff4,
        64'h7593f51f_f0ef0ff5,
        64'hf5930084_559bf5df,
        64'hf0ef0ff5_f5930104,
        64'h559bf69f_f0ef4501,
        64'h0ff5f593_0184559b,
        64'hfee79be3_078500c6,
        64'h802300f1_06b30800,
        64'h0713567d_47810209,
        64'hd993842e_84aae55e,
        64'he95aed56_f152f94a,
        64'he586fd26_e1a20206,
        64'h1993f54e_71558082,
        64'h91411542_8d3d8ff9,
        64'h0057979b_17016709,
        64'h0107d79b_0105179b,
        64'h4105551b_0105151b,
        64'h8d2d00c5_95138da9,
        64'h893d0045_d51b8da9,
        64'h91411542_8d5d0522,
        64'h0085579b_808207f5,
        64'h75138d2d_00451593,
        64'h8d2d8d3d_0045d51b,
        64'h0075d79b_8de98082,
        64'h0141853e_640260a2,
        64'h4781c111_57f5f89f,
        64'hf0efc511_57f9efbf,
        64'hf0efc911_57fdeb7f,
        64'hf0effc6d_e03ff0ef,
        64'h347d4429_b8dff0ef,
        64'hbb050513_00002517,
        64'hc89ff0ef_e022e406,
        64'h11418082_61050015,
        64'h351364a2_644260e2,
        64'h0004051b_fc940ce3,
        64'he37ff0ef_eb3ff0ef,
        64'hbd850513_00002517,
        64'h85aa842a_e53ff0ef,
        64'h02900513_400005b7,
        64'h07700613_fbdff0ef,
        64'h4485e822_ec06e426,
        64'h11018082_01410015,
        64'h3513157d_640260a2,
        64'h0004051b_ef3ff0ef,
        64'hc1250513_85a20000,
        64'h2517e89f_f0ef842a,
        64'he97ff0ef_e022e406,
        64'h03700513_45810650,
        64'h06131141_80826105,
        64'h690264a2_644260e2,
        64'h00153513_f5650513,
        64'h0004051b_01249863,
        64'h88bd00f9_1b634501,
        64'h4785ec9f_f0efecdf,
        64'hf0ef842a_ed3ff0ef,
        64'h84aaed9f_f0efeddf,
        64'hf0efee1f_f0ef892a,
        64'heefff0ef_e04ae426,
        64'he822ec06_45211aa0,
        64'h05930870_06131101,
        64'hbfcd4501_80826105,
        64'h690264a2_644260e2,
        64'h4505f89f_f0ef4585,
        64'hca050513_00002517,
        64'hfe9915e3_c00df25f,
        64'hf0ef892a_347df35f,
        64'hf0ef4501_45810950,
        64'h06134485_71040413,
        64'he04aec06_e4266409,
        64'he8221101_ccdff06f,
        64'h6105c9a5_05130000,
        64'h251760e2_6442da3f,
        64'hf0ef852e_65a2ce7f,
        64'hf0efce25_05130000,
        64'h2517cf3f_f0ef8522,
        64'hcf9ff0ef_e42eec06,
        64'hce850513_00002517,
        64'h842ae822_11018082,
        64'h614564e2_740270a2,
        64'hf47d147d_0007d463,
        64'h4187d79b_0185179b,
        64'hfa7ff0ef_eb5ff0ef,
        64'h85320640_04136622,
        64'hec1ff0ef_0ff47513,
        64'hec9ff0ef_0ff57513,
        64'h0084551b_ed5ff0ef,
        64'h0ff57513_0104551b,
        64'hee1ff0ef_0ff57513,
        64'h0184551b_eedff0ef,
        64'h0404e513_febff0ef,
        64'h84aa842e_ec26f022,
        64'he432f406_7179f07f,
        64'hf06f0ff0_05138082,
        64'h557db7e9_00d70023,
        64'h078500f6_073306c8,
        64'h2683ff79_8b055178,
        64'hbf4dd6b8_07850007,
        64'hc7038082_4501d3b8,
        64'h4719dbb8_577d2000,
        64'h07b700b6_ef630007,
        64'h869b2000_08372000,
        64'h0537fff5_8b85537c,
        64'h20000737_d3b82000,
        64'h07b71060_0713fff5,
        64'h37fd0001_03200793,
        64'h04b76163_40a7873b,
        64'h87aa2000_06b7dbb8,
        64'h57792000_07b706b7,
        64'hec631000_07938082,
        64'h610564a2_d3b84719,
        64'hdbb86442_60e20ff4,
        64'h7513577d_200007b7,
        64'he21ff0ef_dec50513,
        64'h00002517_eafff0ef,
        64'h91011502_4088e37f,
        64'hf0efe0a5_05130000,
        64'h2517e395_8b852401,
        64'h53fc57e0_ff658b05,
        64'h06478493_53f8d3b8,
        64'h10600713_200007b7,
        64'hfff537fd_00010640,
        64'h0793d7a8_dbb85779,
        64'he426e822_ec062000,
        64'h07b71101_e7dff06f,
        64'h6105e3a5_05130000,
        64'h251764a2_60e26442,
        64'hd03c4799_e95ff0ef,
        64'he6050513_00002517,
        64'hf23ff0ef_91010204,
        64'h95132481_eadff0ef,
        64'he5850513_00002517,
        64'h5064d03c_16600793,
        64'hec1ff0ef_e8c50513,
        64'h00002517_f4fff0ef,
        64'h91010204_95132481,
        64'hed9ff0ef_e8450513,
        64'h00002517_5064d03c,
        64'h10400793_20000437,
        64'hfff537fd_000147a9,
        64'hc3b84729_200007b7,
        64'hf01ff0ef_e426e822,
        64'hec06ea45_05131101,
        64'h00002517_80824108,
        64'h8082c10c_ec5ff06f,
        64'h80826105_60e2ecff,
        64'hf0ef0091_4503ed7f,
        64'hf0ef0081_4503f55f,
        64'hf0efec06_002c1101,
        64'h80826145_694264e2,
        64'h740270a2_fe9410e3,
        64'hef9ff0ef_00914503,
        64'hf01ff0ef_34610081,
        64'h4503f81f_f0ef0ff5,
        64'h7513002c_00895533,
        64'h54e10380_0413892a,
        64'hf406e84a_ec26f022,
        64'h71798082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3f3bf_f0ef0091,
        64'h4503f43f_f0ef3461,
        64'h00814503_fc3ff0ef,
        64'h0ff57513_002c0089,
        64'h553b54e1_4461892a,
        64'hf406e84a_ec26f022,
        64'h71798082_00f58023,
        64'h0007c783_00e580a3,
        64'h97aa8111_00074703,
        64'h973e00f5_771326e7,
        64'h87930000_1797b7f5,
        64'h0405f93f_f0ef8082,
        64'h01416402_60a2e509,
        64'h00044503_842ae406,
        64'he0221141_808200e7,
        64'h88230200_071300e7,
        64'h8423fc70_071300e7,
        64'h862300a7_82230ff5,
        64'h751300d7_80230085,
        64'h551b0ff5_769300d7,
        64'h8623f800_06930007,
        64'h822301e7_1793470d,
        64'h02b5553b_0045959b,
        64'h808200a7_8023df65,
        64'h02077713_0147c703,
        64'h07fa478d_80820205,
        64'h75130147_c50307fa,
        64'h478d8082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_100004b7,
        64'h48858593_00001597,
        64'hf1402573_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_372010ef,
        64'h40000137_03249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
