/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 3134;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00000078_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000078_36313025,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000078_36313025,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_78323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000a64_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h00000a64_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_0000000a,
        64'h78363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h0000000a_78363130,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h0000000a_78363130,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_00000a64,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_00000a64,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_00000a64,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_00000a64,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h00000000_00000a78,
        64'h25202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h00000000_0a642520,
        64'h3a737574_61747320,
        64'h2c64656c_69616620,
        64'h64616552_20304453,
        64'h00000000_0a216465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a6425,
        64'h203a7375_74617473,
        64'h202c6465_6c696166,
        64'h206e6f69_74617a69,
        64'h6c616974_696e6920,
        64'h64726163_20304453,
        64'h0000000a_6425203a,
        64'h73757461_7473202c,
        64'h64656c69_6166206c,
        64'h61697469_6e692067,
        64'h69666e6f_63204453,
        64'h00000000_0000000a,
        64'h2164656c_69616620,
        64'h6769666e_6f632070,
        64'h756b6f6f_6c204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_002e2e2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd0080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h08090000_38000000,
        64'hda0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0000a001_fe9fb0ef,
        64'h1a050513_00001517,
        64'h840259a5_85930000,
        64'h05971000_0437e901,
        64'hd82fb0ef_10000537,
        64'h65a180ef_c0ef21e5,
        64'h05130000_151781af,
        64'hc0ef1ca5_05130000,
        64'h1517914f_c0ef2404,
        64'h051382ef_c0ef1de5,
        64'h05130000_1517928f,
        64'hc0ef2404_0513000f,
        64'h4437846f_c0ef1ce5,
        64'h05130000_1517ce0f,
        64'hb0efe022_e406a005,
        64'h05132005_85931141,
        64'h02626537_65f18082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'h96afc0ef_4505a031,
        64'hfef42623_4785e789,
        64'h27810807_f7932781,
        64'h87aaa31f_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h37830001_a011f6e7,
        64'hfee30270_07930ff7,
        64'hf713fe94_4783fef4,
        64'h04a32785_fe944783,
        64'hcf992781_0407f793,
        64'h278187aa_a6bfe0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_a0adfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaa61f_d0effd84,
        64'h35035007_85936785,
        64'h46014685_a829fef4,
        64'h262387aa_a7bfd0ef,
        64'hfd843503_30078593,
        64'h67854601_468500f7,
        64'h1f634785_873e0347,
        64'hc783fd84_3783a8ad,
        64'hfe0404a3_a26fc0ef,
        64'h4505b13f_e0ef853e,
        64'h03e00593_863afe64,
        64'h570343dc_fd843783,
        64'hfef41323_0407e793,
        64'hfe645783_fef41323,
        64'h87aab01f_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h378366e7_92234741,
        64'h00000797_b55fe0ef,
        64'h853e4591_863afea4,
        64'h570343dc_fd843783,
        64'hfef41523_8ff917fd,
        64'h6785fea4_5703fef4,
        64'h15230017_979bfea4,
        64'h5783aa35_478568e7,
        64'hae234705_00000797,
        64'h9bcfc0ef_74c50513,
        64'h00000517_74458593,
        64'h00000597_48e00613,
        64'ha02502f7_1c63478d,
        64'h873e0377_c783fd84,
        64'h3783fef4_15230400,
        64'h07936c07_ab230000,
        64'h0797a251_47856ee7,
        64'ha2234705_00000797,
        64'ha04fc0ef_79450513,
        64'h00000517_78c58593,
        64'h00000597_48d00613,
        64'ha02504f7_17631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_37837007,
        64'had230000_0797c385,
        64'hfd843783_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aab8ff_e0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783c4ff,
        64'he0ef853e_03000593,
        64'h460943dc_fd843783,
        64'hdfc52781_8b89fe84,
        64'h2783a83d_fef42623,
        64'h4785c73f_e0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hc3852781_8ff967a1,
        64'hfe842703_fef42423,
        64'h87aac61f_e0ef853e,
        64'h03000593_43dcfd84,
        64'h3783a8bd_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hc57fd0ef_fd843503,
        64'h60000593_863e4681,
        64'hfd442783_fcf42a23,
        64'h87aefca4_3c231800,
        64'hf022f406_71798082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'hc55fe0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfc843783_d15fe0ef,
        64'h853e0300_05934609,
        64'h43dcfc84_3783dfc5,
        64'h27818b89_fdc42783,
        64'ha83dfef4_26234785,
        64'hd39fe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fc84_3783c385,
        64'h27818ff9_67a1fdc4,
        64'h2703fcf4_2e2387aa,
        64'hd27fe0ef_853e0300,
        64'h059343dc_fc843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aad1df,
        64'hd0effc84_35038007,
        64'h85936785_863e4685,
        64'hfe442783_8ae79b23,
        64'h47450000_1797f56f,
        64'he0effc84_350385be,
        64'hfc043603_2781fe24,
        64'h5783dbbf_e0ef853e,
        64'h4591863a_fe045703,
        64'h43dcfc84_3783fef4,
        64'h10238ff9_17fd6785,
        64'hfe045703_fef41023,
        64'h20000793_fef41123,
        64'h4785fce7_dee31ff0,
        64'h07930007_871bfe84,
        64'h2783fef4_24232785,
        64'hfe842783_00078023,
        64'h97bafc04_3703fe84,
        64'h2783a215_478592e7,
        64'ha6234705_00001797,
        64'hc4cfc0ef_9dc50513,
        64'h00001517_9d458593,
        64'h00001597_35d00613,
        64'ha081fe04_24239407,
        64'ha9230000_1797aaa1,
        64'h478596e7_a0234705,
        64'h00001797_c80fc0ef,
        64'ha1050513_00001517,
        64'ha0858593_00001597,
        64'h35c00613_a02502f7,
        64'h1d631117_87931111,
        64'h17b7873e_53dcfc84,
        64'h37839807_ab230000,
        64'h1797c385_fc843783,
        64'hfe042223_fcb43023,
        64'hfca43423_0080f822,
        64'hfc067139_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623a019,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_e63fd0ef,
        64'hfd843503_a0078593,
        64'h67ad4601_4681a03d,
        64'hfef42623_4785a82d,
        64'h4785a0e7_a0234705,
        64'h00001797_d20fc0ef,
        64'hab050513_00001517,
        64'haa858593_00001597,
        64'h32d00613_a025cb8d,
        64'h2781fec4_2783fef4,
        64'h262387aa_eb3fd0ef,
        64'hfd843503_70078593,
        64'h678d863e_46814bbc,
        64'hfd843783_a407a423,
        64'h00001797_a8414785,
        64'ha4e7ab23_47050000,
        64'h1797d76f_c0efb065,
        64'h05130000_1517afe5,
        64'h85930000_159732c0,
        64'h0613a025_04f71e63,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'ha807a623_00001797,
        64'hc385fd84_3783fca4,
        64'h3c231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_fe842783,
        64'hfe042423_fa5fe0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0047e793,
        64'hfe445783_43d8fd84,
        64'h3783fef4_122387aa,
        64'hf8ffe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'hd3e52781_8b892781,
        64'hfe645783_fef41323,
        64'h87aafb1f_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783a821_fef41323,
        64'h87aafc9f_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783812f_f0ef853e,
        64'h02c00593_863afe44,
        64'h570343dc_fd843783,
        64'hfef41223_0017e793,
        64'h93c117c2_8fd9fe44,
        64'h5783fec4_5703fef4,
        64'h1623f007_f793fec4,
        64'h5783fef4_16230087,
        64'h979bfec4_5783fef4,
        64'h12230ff7_f793fe44,
        64'h5783fef4_122387aa,
        64'h82eff0ef_853e02c0,
        64'h059343dc_fd843783,
        64'ha0a587af_f0ef853e,
        64'h02c00593_863afe44,
        64'h570343dc_fd843783,
        64'hfef41223_0017e793,
        64'h93c117c2_8fd9fe44,
        64'h57839341_03079713,
        64'h8fd9fe24_5783fec4,
        64'h5703fef4_1623f007,
        64'hf793fec4_5783fef4,
        64'h16230087_979bfec4,
        64'h5783fef4_11230c07,
        64'hf793fe24_5783fef4,
        64'h11230067_979bfe24,
        64'h5783fef4_11230087,
        64'hd79bfec4_5783fef4,
        64'h122303f7_f793fe44,
        64'h5783fef4_122387aa,
        64'h8c6ff0ef_853e02c0,
        64'h059343dc_fd843783,
        64'h08f71e63_4789873e,
        64'h0367c783_fd843783,
        64'ha249fef4_24234785,
        64'h00e7f663_10000793,
        64'h0007871b_fee45783,
        64'hfae7fee3_10000793,
        64'h0007871b_fee45783,
        64'hfef41723_0017979b,
        64'hfee45783_a839fef4,
        64'h16230017_d79bfee4,
        64'h578300e7_e9632781,
        64'hfd442783_0007871b,
        64'h02f757bb_2781fee4,
        64'h57834798_fd843783,
        64'ha82dfef4_17234785,
        64'ha2edfef4_24234785,
        64'h06e7fa63_7fe00793,
        64'h0007871b_fee45783,
        64'hfae7ffe3_7fe00793,
        64'h0007871b_fee45783,
        64'hfef41723_2785fee4,
        64'h5783a831_fef41623,
        64'h0017d79b_fee45783,
        64'h00e7e963_2781fd44,
        64'h27830007_871b02f7,
        64'h57bb2781_fee45783,
        64'h4798fd84_3783a825,
        64'hfef41723_4785ac91,
        64'h4785d0e7_a4234705,
        64'h00001797_829fc0ef,
        64'hdb850513_00001517,
        64'hdb058593_00001597,
        64'h2b800613_a02508f7,
        64'h19634789_873e0367,
        64'hc783fd84_3783a26f,
        64'hf0ef853e_02c00593,
        64'h863afe44_570343dc,
        64'hfd843783_fef41223,
        64'h9be9fe44_5783fef4,
        64'h122387aa_a12ff0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_d607a823,
        64'h00001797_a4e94785,
        64'hd6e7af23_47050000,
        64'h179789ff_c0efe2e5,
        64'h05130000_1517e265,
        64'h85930000_15972b70,
        64'h0613a025_06f71e63,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'hda07aa23_00001797,
        64'hc385fd84_3783fe04,
        64'h1623fcf4_2a2387ae,
        64'hfca43c23_1800f022,
        64'hf4067179_80826165,
        64'h740670a6_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aaa32f,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcf984,
        64'h3783b72f_f0ef853e,
        64'h02800593_863a0ff7,
        64'h7713fe44_270343dc,
        64'hf9843783_fef42223,
        64'h0047e793_fe442783,
        64'hfef42223_87aab64f,
        64'hf0ef853e_02800593,
        64'h43dcf984_3783a49f,
        64'hc0ef3e80_0513a09d,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_730000ef,
        64'hf9843503_02f71163,
        64'h479d873e_57fcf984,
        64'h3783a849_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h0b8000ef_f9843503,
        64'h85be5f9c_f9843783,
        64'hb88ff0ef_853e0300,
        64'h05934609_43dcf984,
        64'h3783dfc5_27818b89,
        64'hfe442783_a8d1fef4,
        64'h26234785_bacff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8f984,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_b9aff0ef,
        64'h853e0300_059343dc,
        64'hf9843783_aa11fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aab90f_e0eff984,
        64'h35036000_0593863e,
        64'h4681fe84_2783df98,
        64'h5007071b_03197737,
        64'hf9843783_fef42423,
        64'h1007879b_03b907b7,
        64'ha831df98_5007071b,
        64'h03197737_f9843783,
        64'hfef42423_1007879b,
        64'h03b907b7_02f71063,
        64'h4791873e_57fcf984,
        64'h3783a099_df982007,
        64'h071b0beb_c737f984,
        64'h3783fef4_24232007,
        64'h879b03b9_07b702f7,
        64'h1063479d_873e57fc,
        64'hf9843783_a275fef4,
        64'h26234785_14078963,
        64'h2781fec4_2783fef4,
        64'h262387aa_1d4000ef,
        64'hf9843503_50078593,
        64'h031977b7_df985007,
        64'h071b0319_7737f984,
        64'h3783cb2f_f0ef853e,
        64'h03000593_460943dc,
        64'hf9843783_dfc52781,
        64'h8b89fe44_2783aafd,
        64'hfef42623_4785cd6f,
        64'hf0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hf9843783_c3852781,
        64'h8ff967a1_fe442703,
        64'hfef42223_87aacc4f,
        64'hf0ef853e_03000593,
        64'h43dcf984_3783ac3d,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_cbafe0ef,
        64'hf9843503_60000593,
        64'h863e4681_fe842783,
        64'hfef42423_1007879b,
        64'h03b907b7_0cf71663,
        64'h4789873e_0347c783,
        64'hf9843783_a451fef4,
        64'h26234785_22078563,
        64'h2781fec4_2783fef4,
        64'h262387aa_2ac000ef,
        64'hf9843503_85be5f9c,
        64'hf9843783_df980807,
        64'h071b02fa_f737f984,
        64'h3783d8af_f0ef853e,
        64'h03000593_460943dc,
        64'hf9843783_dfc52781,
        64'h8b89fe44_2783acd9,
        64'hfef42623_4785daef,
        64'hf0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hf9843783_c3852781,
        64'h8ff967a1_fe442703,
        64'hfef42223_87aad9cf,
        64'hf0ef853e_03000593,
        64'h43dcf984_3783ae19,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_d92fe0ef,
        64'hf9843503_60000593,
        64'h863e4685_fe842783,
        64'hfef42423_37c58100,
        64'h07b712e7_9a234745,
        64'h00001797_fd5fe0ef,
        64'hf9843503_85be863a,
        64'hfa040713_2781fe24,
        64'h5783e3af_f0ef853e,
        64'h4591863a_fe045703,
        64'h43dcf984_3783fef4,
        64'h10238ff9_17fd6785,
        64'hfe045703_fef41023,
        64'h04000793_fef41123,
        64'h4785ae79_478518e7,
        64'ha2234705_00001797,
        64'hca5fc0ef_23450513,
        64'h00001517_22c58593,
        64'h00001597_1f400613,
        64'ha02514f7_11634785,
        64'h873e0347_c783f984,
        64'h37831a07_ab230000,
        64'h1797aef9_47851ce7,
        64'ha2234705_00001797,
        64'hce5fc0ef_27450513,
        64'h00001517_26c58593,
        64'h00001597_1f300613,
        64'ha02504f7_13631117,
        64'h87931111_17b7873e,
        64'h53dcf984_37831e07,
        64'had230000_1797c385,
        64'hf9843783_fc043c23,
        64'hfc043823_fc043423,
        64'hfc043023_fa043c23,
        64'hfa043823_fa043423,
        64'hfa043023_f8a43c23,
        64'h1880f0a2_f4867159,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aae8ef_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfc84_3783f4ef,
        64'hf0ef853e_03000593,
        64'h460943dc_fc843783,
        64'hdfc52781_8b89fdc4,
        64'h2783a83d_fef42623,
        64'h4785f72f_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fc843783,
        64'hc3852781_8ff967a1,
        64'hfdc42703_fcf42e23,
        64'h87aaf60f_f0ef853e,
        64'h03000593_43dcfc84,
        64'h3783a8bd_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hf56fe0ef_fc843503,
        64'h60000593_863e4685,
        64'hfe042783_fef42023,
        64'h37c10100_07b72ee7,
        64'h9c234745_00001797,
        64'h998ff0ef_fc843503,
        64'h85befc04_36032781,
        64'hfe645783_ffcff0ef,
        64'h853e4591_863afe44,
        64'h570343dc_fc843783,
        64'hfef41223_8ff917fd,
        64'h6785fe44_5703fef4,
        64'h12230400_0793fef4,
        64'h13234785_fce7dee3,
        64'h03f00793_0007871b,
        64'hfe842783_fef42423,
        64'h2785fe84_27830007,
        64'h802397ba_fc043703,
        64'hfe842783_a2354785,
        64'h36e7a723_47050000,
        64'h1797e8ff_c0ef41e5,
        64'h05130000_15174165,
        64'h85930000_15971a00,
        64'h0613a081_fe042423,
        64'h3807aa23_00001797,
        64'ha2854785_3ae7a123,
        64'h47050000_1797ec3f,
        64'hc0ef4525_05130000,
        64'h151744a5_85930000,
        64'h159719f0_0613a025,
        64'h02f71d63_11178793,
        64'h111117b7_873e53dc,
        64'hfc843783_3c07ac23,
        64'h00001797_c385fc84,
        64'h3783fcb4_3023fca4,
        64'h34230080_f822fc06,
        64'h71398082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_851ff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fd843783,
        64'h911ff0ef_853e03e0,
        64'h0593863a_93411742,
        64'hfe842703_43dcfd84,
        64'h3783fef4_24238fd9,
        64'hfe842783_57f8fd84,
        64'h3783fef4_24238ff9,
        64'h17e167c1_fe842703,
        64'hfef42423_87aa915f,
        64'hf0ef853e_03e00593,
        64'h43dcfd84_378304f7,
        64'h19634791_873e57fc,
        64'hfd843783_9edff0ef,
        64'h853e0280_0593863a,
        64'h0ff77713_fe842703,
        64'h43dcfd84_3783fef4,
        64'h24230027_e793fe84,
        64'h2783a039_fef42423,
        64'h0207e793_fe842783,
        64'h00f71963_478d873e,
        64'h0377c783_fd843783,
        64'hfef42423_87aa9fdf,
        64'hf0ef853e_02800593,
        64'h43dcfd84_37838e0f,
        64'hd0ef3e80_05139cff,
        64'hf0ef853e_03000593,
        64'h460943dc_fd843783,
        64'hdfc52781_8b89fe84,
        64'h2783a8f5_fef42623,
        64'h47859f3f_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hc3852781_8ff967a1,
        64'hfe842703_fef42423,
        64'h87aa9e1f_f0ef853e,
        64'h03000593_43dcfd84,
        64'h3783aa35_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h9d7fe0ef_fd843503,
        64'h60000593_863e4681,
        64'hfe442783_fef42223,
        64'h1007879b_03b707b7,
        64'ha039fef4_22235007,
        64'h879b03b7_07b700f7,
        64'h19634791_873e57fc,
        64'hfd843783_a02dfef4,
        64'h22232007_879b03b7,
        64'h07b7a825_fef42223,
        64'h6007879b_03b707b7,
        64'h00f71963_4791873e,
        64'h57fcfd84_378302f7,
        64'h1763478d_873e0377,
        64'hc783fd84_378302e7,
        64'h8ba34709_fd843783,
        64'ha03102e7_8ba3470d,
        64'hfd843783_00f71863,
        64'h47a1873e_4bdcfd84,
        64'h378300f7_1f634795,
        64'h873e0347_c783fd84,
        64'h378302f7_17634789,
        64'h873e0367_c783fd84,
        64'h3783a431_fef42623,
        64'h47851207_8c632781,
        64'hfec42783_fef42623,
        64'h87aaaa9f_e0effd84,
        64'h35036007_859367a1,
        64'h863e4681_fe442783,
        64'hfef42223_0377c783,
        64'hfd843783_02e78ba3,
        64'h4709fd84_3783ac81,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_aebfe0ef,
        64'hfd843503_70078593,
        64'h678d863e_46814bbc,
        64'hfd843783_06f71b63,
        64'h4785873e_0347c783,
        64'hfd843783_a479fe04,
        64'h262300e7_e563478d,
        64'h873e4bdc_fd843783,
        64'ha45d4785_6ae7a523,
        64'h47050000_17979caf,
        64'hd0ef75a5_05130000,
        64'h15177525_85930000,
        64'h15971130_0613a025,
        64'h04f71063_4789873e,
        64'h0367c783_fd843783,
        64'h6c07ae23_00001797,
        64'ha4dd4785_6ee7a523,
        64'h47050000_1797a0af,
        64'hd0ef79a5_05130000,
        64'h15177925_85930000,
        64'h15971120_0613a025,
        64'h04f71363_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_7207a023,
        64'h00001797_c385fd84,
        64'h3783fca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'hb95ff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_c55ff0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe042783,
        64'ha83dfef4_26234785,
        64'hc79ff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe04,
        64'h2703fef4_202387aa,
        64'hc67ff0ef_853e0300,
        64'h059343dc_fd843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aac5df,
        64'he0effd84_35033007,
        64'h859367ad_460186be,
        64'h2781fe64_57837ee7,
        64'h9c234745_00001797,
        64'he98ff0ef_fd843503,
        64'h85befd04_36032781,
        64'hfe645783_cfdff0ef,
        64'h853e4591_863afe44,
        64'h570343dc_fd843783,
        64'hfef41223_8ff917fd,
        64'h6785fe44_5703fef4,
        64'h122347a1_fef41323,
        64'h4785a8e5_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hcd7fe0ef_fd843503,
        64'h70078593_678d863e,
        64'h46814bbc_fd843783,
        64'hfce7dfe3_479d0007,
        64'h871bfe84_2783fef4,
        64'h24232785_fe842783,
        64'h00078023_97bafd04,
        64'h3703fe84_2783aa81,
        64'h478588e7_ac234705,
        64'h00002797_bb8fd0ef,
        64'h94850513_00002517,
        64'h94058593_00002597,
        64'h0ba00613_a081fe04,
        64'h24238a07_af230000,
        64'h2797a251_47858ce7,
        64'ha6234705_00002797,
        64'hbecfd0ef_97c50513,
        64'h00002517_97458593,
        64'h00002597_0b900613,
        64'ha02502f7_1d631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_37839007,
        64'ha1230000_2797c385,
        64'hfd843783_fcb43823,
        64'hfca43c23_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623e1ff,
        64'hf0ef8536_4591863e,
        64'h93c117c2_8ff917fd,
        64'h6785fd64_570343d4,
        64'hfd843783_fef42623,
        64'h278187aa_d99ff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fd843783,
        64'ha081fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aae05f,
        64'he0effd84_35036585,
        64'h863e4681_2781fd64,
        64'h5783a0ad_fef42623,
        64'h4785a89d_47859ae7,
        64'ha2234705_00002797,
        64'hcc4fd0ef_a5450513,
        64'h00002517_a4c58593,
        64'h00002597_07f00613,
        64'ha025cb8d_27813037,
        64'hf793fe84_2783fef4,
        64'h242387aa_e19ff0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h37839e07_a7230000,
        64'h2797a0f9_47859ee7,
        64'hae234705_00002797,
        64'hd1cfd0ef_aac50513,
        64'h00002517_aa458593,
        64'h00002597_07e00613,
        64'ha02504f7_1f631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783a207,
        64'ha9230000_2797c385,
        64'hfd843783_fcf41b23,
        64'h87aefca4_3c231800,
        64'hf022f406_71798082,
        64'h61056442_60e20001,
        64'heb7ff0ef_853e85ba,
        64'hfea44703_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h052387ba_fef405a3,
        64'h87b6fef4_26238732,
        64'h86ae87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_853e87aa,
        64'hea9ff0ef_853e9381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef405a3_87bafef4,
        64'h2623872e_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e20001,
        64'hf63ff0ef_853e85ba,
        64'hfe845703_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h142387ba_fef405a3,
        64'h87b6fef4_26238732,
        64'h86ae87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_853e87aa,
        64'hf47ff0ef_853e9381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef405a3_87bafef4,
        64'h2623872e_87aa1000,
        64'he822ec06_11018082,
        64'h61457422_000100e7,
        64'h9023fd64_5703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_1b2387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61457422,
        64'h000100e7_8023fd74,
        64'h4703fe84_3783fef4,
        64'h3423fd84_3783fcf4,
        64'h0ba387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61056462_853e2781,
        64'h439cfe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826105_6462853e,
        64'h93c117c2_0007d783,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61056462_853e0ff7,
        64'hf7930007_c783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826161,
        64'h640660a6_853efec4,
        64'h2783fe04_2623d3f8,
        64'hfb843783_0007871b,
        64'h0097d79b_fd842783,
        64'hfcf42c23_02f707bb,
        64'hfe042783_fd842703,
        64'hfcf42c23_02f707bb,
        64'hfdc42703_27812785,
        64'hfd842783_fcf42c23,
        64'h8fd9fd84_27830007,
        64'h871b8ff9_c0078793,
        64'h6785873e_278100a7,
        64'h979bfd04_2783fcf4,
        64'h2c230167_d79bfcc4,
        64'h2783fcf4_2e232781,
        64'h00f717bb_47052781,
        64'h27892781_8b9d2781,
        64'h0077d79b_fcc42783,
        64'hfef42023_278100f7,
        64'h17bb4705_27818bbd,
        64'h27810087_d79bfd04,
        64'h278302e7_8aa3fb84,
        64'h37830ff7_f7138bbd,
        64'h0ff7f793_27810127,
        64'hd79bfd44_2783fcf4,
        64'h2a232781_87aa9bdf,
        64'hd0ef853e_93811782,
        64'h278127f1_43dcfb84,
        64'h3783fcf4_28232781,
        64'h87aa9d9f_d0ef853e,
        64'h93811782_278127e1,
        64'h43dcfb84_3783fcf4,
        64'h26232781_87aa9f5f,
        64'hd0ef853e_93811782,
        64'h278127d1_43dcfb84,
        64'h3783fcf4_24232781,
        64'h87aaa11f_d0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783a23d,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_9d2ff0ef,
        64'hfb843503_90078593,
        64'h6785863e_46814bbc,
        64'hfb843783_aab1fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaa00f_f0effb84,
        64'h35033000_0593863e,
        64'h46814bbc_fb843783,
        64'hcbb81234_0737fb84,
        64'h3783c7f8_fb843783,
        64'h0007871b_87aab31f,
        64'hd0ef853e_45f143dc,
        64'hfb843783_c7b8fb84,
        64'h37830007_871b87aa,
        64'hb4bfd0ef_853e45e1,
        64'h43dcfb84_3783c3f8,
        64'hfb843783_0007871b,
        64'h87aab65f_d0ef853e,
        64'h45d143dc_fb843783,
        64'hc3b8fb84_37830007,
        64'h871b87aa_b7ffd0ef,
        64'h853e45c1_43dcfb84,
        64'h3783aaed_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'ha9eff0ef_fb843503,
        64'h20000593_46014681,
        64'hdb984705_fb843783,
        64'hc7892781_8ff94000,
        64'h07b7fe84_2703fa07,
        64'hdde3fe84_2783fef4,
        64'h242387aa_b3bfd0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'haca1fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaafcf,
        64'hf0effb84_35031000,
        64'h059340ff_86374681,
        64'ha091fe04_2423a459,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_b2aff0ef,
        64'hfb843503_45814601,
        64'h4681a46d_fef42623,
        64'h4785e789_27818ff9,
        64'h67c1fe44_2703fef4,
        64'h222387aa_bbbfd0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfb84,
        64'h3783cb8d_47dcfb84,
        64'h378302f7_0e634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfb843783_a6014785,
        64'hf0e7a723_47050000,
        64'h2797a2ff_d0eff9e5,
        64'h05130000_2517f9e5,
        64'h85930000_25976710,
        64'h0613a025_04f71363,
        64'h4789873e_0367c783,
        64'hfb843783_f407a023,
        64'h00002797_a6814785,
        64'hf4e7a723_47050000,
        64'h2797a6ff_d0effde5,
        64'h05130000_2517fde5,
        64'h85930000_25976700,
        64'h0613a025_04f71363,
        64'h11178793_111117b7,
        64'h873e53dc_fb843783,
        64'hf807a223_00002797,
        64'hc385fb84_3783faa4,
        64'h3c230880_e0a2e486,
        64'h715d8082_61217442,
        64'h70e20001_d05fd0ef,
        64'h853a85be_27810807,
        64'h8793fd84_37839301,
        64'h02079713_27810587,
        64'h879b43dc_fd843783,
        64'h00e79123_97b6078e,
        64'h07c19381_02061793,
        64'hfd843683_93410307,
        64'h971302f7_07bb0006,
        64'h861b36fd_fec42683,
        64'h93c117c2_fe442783,
        64'h93410307_9713fd44,
        64'h278300e7_90230230,
        64'h071397ba_078e07c1,
        64'h93811782_fd843703,
        64'h278137fd_fec42783,
        64'hc3d897b6_078e07c1,
        64'h93810206_1793fd84,
        64'h36830007_871b9fb9,
        64'h0006861b_36fdfec4,
        64'h26832781_0107979b,
        64'hfe842783_0007871b,
        64'hfc843783_f8e7ebe3,
        64'h2781fe84_27830007,
        64'h871b37fd_fec42783,
        64'hfef42423_2785fe84,
        64'h27830007_912397ba,
        64'h078e07c1_fe846783,
        64'hfd843703_00e79023,
        64'h02100713_97ba078e,
        64'h07c1fe84_6783fd84,
        64'h3703c3d8_97b6078e,
        64'h07c1fe84_6783fd84,
        64'h36830007_871b9fb9,
        64'h27810107_979bfe84,
        64'h27830007_871bfc84,
        64'h3783a8b1_fe042423,
        64'hfef42623_2785fec4,
        64'h2783c791_27818ff9,
        64'h17fd67c1_873e2781,
        64'h02f707bb_fe442783,
        64'hfd442703_fef42623,
        64'h0107d79b_278102f7,
        64'h07bbfe44_2783fd44,
        64'h2703a835_fef42623,
        64'h478500f7_766367c1,
        64'h873e2781_02f707bb,
        64'hfe442783_fd442703,
        64'hfef42223_8ff917fd,
        64'h6785fe44_2703fef4,
        64'h222387aa_ebffd0ef,
        64'h853e4591_43dcfd84,
        64'h3783fe04_2223fe04,
        64'h2423fe04_2623fcf4,
        64'h2a23fcc4_342387ae,
        64'hfca43c23_0080f822,
        64'hfc067139_80826145,
        64'h740270a2_853efec4,
        64'h27830001_a011fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aae10f_f0effd84,
        64'h35037000_0593863e,
        64'h46814bbc_fd843783,
        64'hfe042623_fca43c23,
        64'h1800f022_f4067179,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623f87f_d0ef853e,
        64'h03000593_460943dc,
        64'hfd843783_dfc52781,
        64'h8b89fe44_2783a00d,
        64'hfef42623_4785fabf,
        64'hd0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c3852781,
        64'h8ff967a1_fe442703,
        64'hfef42223_87aaf99f,
        64'hd0ef853e_03000593,
        64'h43dcfd84_3783a08d,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_ebaff0ef,
        64'hfd843503_90078593,
        64'h6789863e_86bafd44,
        64'h2783fd04_270324e7,
        64'h9d230270_07130000,
        64'h2797a879_fef42623,
        64'h4785c3b9_2781fec4,
        64'h2783fef4_262387aa,
        64'hef6ff0ef_fd843503,
        64'h80078593_6789863e,
        64'h86bafd44_2783fd04,
        64'h270328e7_9a23470d,
        64'h00002797_02f71f63,
        64'h47850007_871bfd04,
        64'h27831420_00effd84,
        64'h350385be_fc843603,
        64'hfd042783_a8e5fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa0810_00effd84,
        64'h35032000_059302f7,
        64'h03632000_0793873e,
        64'h278187aa_fd3fd0ef,
        64'h853e9381_17822781,
        64'h279143dc_fd843783,
        64'haa35fef4_26234785,
        64'he7892781_8ff967c1,
        64'hfe842703_fef42423,
        64'h87aa800f_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'hcb8d47dc_fd843783,
        64'h02f70e63_400007b7,
        64'h873e2781_8ff9c000,
        64'h07b7873e_579cfd84,
        64'h378300f7_1f634789,
        64'h873e0367_c783fd84,
        64'h3783fcf4_282387ba,
        64'hfcf42a23_fcd43423,
        64'h873287ae_fca43c23,
        64'h0080f822_fc067139,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aa880f_e0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_378396af,
        64'he0ef853e_03000593,
        64'h460943dc_fd843783,
        64'hdfc52781_8b89fe44,
        64'h2783a83d_fef42623,
        64'h478598ef_e0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aa97cf_e0ef853e,
        64'h03000593_43dcfd84,
        64'h3783a8bd_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h89fff0ef_fd843503,
        64'h20078593_6785863e,
        64'h86bafd44_2783fd04,
        64'h270342e7_9f230370,
        64'h07130000_2797a86d,
        64'hfef42623_4785c3b9,
        64'h2781fec4_2783fef4,
        64'h262387aa_8dbff0ef,
        64'hfd843503_10078593,
        64'h6785863e_86bafd44,
        64'h2783fd04_270346e7,
        64'h9c23474d_00002797,
        64'h02f71f63_47850007,
        64'h871bfd04_27833260,
        64'h00effd84_350385be,
        64'hfc843603_fd042783,
        64'haa11fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa2650,
        64'h00effd84_35032000,
        64'h059302f7_03632000,
        64'h0793873e_278187aa,
        64'h9b6fe0ef_853e9381,
        64'h17822781_279143dc,
        64'hfd843783_aaa1fef4,
        64'h26234785_e7892781,
        64'h8ff967c1_fe842703,
        64'hfef42423_87aa9e4f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_cb8d47dc,
        64'hfd843783_02f70e63,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cfd84_378300f7,
        64'h1f634789_873e0367,
        64'hc783fd84_3783fcf4,
        64'h282387ba_fcf42a23,
        64'hfcd43423_873287ae,
        64'hfca43c23_0080f822,
        64'hfc067139_80826145,
        64'h7422853e_fec42783,
        64'h0001a011_0001a021,
        64'h0001a031_fef42623,
        64'h8fd9fd44_2783fec4,
        64'h2703a831_fef42623,
        64'h01a7e793_fec42783,
        64'ha02dfef4_262303a7,
        64'he793fec4_2783a825,
        64'hfef42623_01a7e793,
        64'hfec42783_a099fef4,
        64'h26230027_e793fec4,
        64'h2783a891_fef42623,
        64'h03a7e793_fec42783,
        64'ha08dfef4_262303a7,
        64'he793fec4_2783a885,
        64'hfef42623_01a7e793,
        64'hfec42783_a8bdfef4,
        64'h26230097_e793fec4,
        64'h2783a071_fef42623,
        64'h03a7e793_fec42783,
        64'ha869fef4_262301a7,
        64'he793fec4_278300f7,
        64'h19634785_873e0347,
        64'hc783fd84_3783a865,
        64'hfef42623_01a7e793,
        64'hfec42783_a0d9fef4,
        64'h262301a7_e793fec4,
        64'h2783a8d1_fef42623,
        64'h01b7e793_fec42783,
        64'ha0cdfef4_262303a7,
        64'he793fec4_278300f7,
        64'h19634785_873e0347,
        64'hc783fd84_3783a201,
        64'hfef42623_01b7e793,
        64'hfec42783_a239fef4,
        64'h262301b7_e793fec4,
        64'h2783aa31_fef42623,
        64'h0097e793_fec42783,
        64'ha22dfef4_26230027,
        64'he793fec4_2783aa39,
        64'h0ef70563_90078793,
        64'h67ad0007_871b10e6,
        64'h8a633007_0713672d,
        64'h0007869b_10e68a63,
        64'ha0070713_672d0007,
        64'h869ba2a9_16f70363,
        64'ha0078793_67910007,
        64'h871b0ee6_8d63d007,
        64'h07136725_0007869b,
        64'h0ae68963_60070713,
        64'h67210007_869b02d7,
        64'h68637007_07136725,
        64'h0007869b_14e68063,
        64'h70070713_67250007,
        64'h869baa49_14f70863,
        64'h80078793_67890007,
        64'h871b18e6_8b634007,
        64'h0713670d_0007869b,
        64'h16e68663_90070713,
        64'h67090007_869baa7d,
        64'h16f70763_20078793,
        64'h67850007_871b16e6,
        64'h8e635007_07136705,
        64'h0007869b_18e68563,
        64'h30070713_67050007,
        64'h869b02d7_68637007,
        64'h07136705_0007869b,
        64'h1ae68a63_70070713,
        64'h67050007_869b06d7,
        64'h6c637007_0713670d,
        64'h0007869b_20e68463,
        64'h70070713_670d0007,
        64'h869ba40d_1cf70263,
        64'hb0078793_67850007,
        64'h871b1ce6_89636705,
        64'h0007869b_1ce68e63,
        64'hc0070713_67050007,
        64'h869ba4a9_1af70263,
        64'h70000793_0007871b,
        64'h1ee68563_90070713,
        64'h67050007_869b1c07,
        64'h06632701_8007871b,
        64'h02d76563_a0070713,
        64'h67050007_869b20e6,
        64'h8f63a007_07136705,
        64'h0007869b_a47118f7,
        64'h08633000_07930007,
        64'h871b1ae6_85635000,
        64'h07130007_869b2ae6,
        64'h8e634000_07130007,
        64'h869bac4d_18f70d63,
        64'h10000793_0007871b,
        64'h2c070963_0007871b,
        64'h00d76d63_20000713,
        64'h0007869b_1ce68463,
        64'h20000713_0007869b,
        64'h04d76c63_60000713,
        64'h0007869b_20e68563,
        64'h60000713_0007869b,
        64'h0cd76d63_10070713,
        64'h67050007_869b2ae6,
        64'h8a631007_07136705,
        64'h0007869b_fd442783,
        64'hfef42623_fd442783,
        64'hfcf42a23_87aefca4,
        64'h3c231800_f4227179,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623e86f_e0ef853e,
        64'h03000593_460543dc,
        64'hfd843783_d3a92781,
        64'h8b85fe04_2783a00d,
        64'hea4fe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783fef4,
        64'h26234789_e7812781,
        64'h9bf9fec4_2783fef4,
        64'h262387aa_e96fe0ef,
        64'h853e0320_059343dc,
        64'hfd843783_c3a12781,
        64'h8ff967a1_fe042703,
        64'ha899eeef_e0ef853e,
        64'h03000593_02000613,
        64'h43dcfd84_3783cf81,
        64'h27810207_f7932781,
        64'h87aaed4f_e0ef853e,
        64'h03000593_43dcfd84,
        64'h378302f7_1b633007,
        64'h87936785_0007871b,
        64'hfd442783_00f70b63,
        64'h50078793_67850007,
        64'h871bfd44_2783fef4,
        64'h202387aa_f0efe0ef,
        64'h853e0300_059343dc,
        64'hfd843783_ef4fe0ef,
        64'h853a85be_27818fd5,
        64'h27819aa7_d7830000,
        64'h37970007_869b0107,
        64'h979bfe44_27839301,
        64'h02079713_278127b1,
        64'h43dcfd84_3783a229,
        64'hfef42623_4785c789,
        64'h27810207_f793fe44,
        64'h2783cb99_27818b89,
        64'hfe842783_fef42423,
        64'h87aaed8f_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'h02f70f63_30078793,
        64'h67850007_871bfd44,
        64'h278304f7_08635007,
        64'h87936785_0007871b,
        64'hfd442783_fef42223,
        64'h8ff917fd_6791fe44,
        64'h2703fef4_222387aa,
        64'h18c000ef_fd843503,
        64'h85befd44_278380bf,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_821fe0ef,
        64'h853a0300_0593fff7,
        64'h861367c1_43d8fd84,
        64'h3783fd2f_e0ef853e,
        64'h85bafd04_27039381,
        64'h17822781_27a143dc,
        64'hfd843783_8d1fe0ef,
        64'h853e02e0_05934639,
        64'h43dcfd84_3783863f,
        64'he0ef853e_4599863a,
        64'h93411742_fcc42703,
        64'h43dcfd84_3783aaed,
        64'hfef42623_4785a419,
        64'h4785ace7_a4234705,
        64'h00003797_de8fe0ef,
        64'hb5850513_00003517,
        64'hb5858593_00003597,
        64'h44c00613_a025cb8d,
        64'h27818b85_fe842783,
        64'hfef42423_87aafe4f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_b007a823,
        64'h00003797_acb14785,
        64'hb0e7af23_47050000,
        64'h3797e3ef_e0efbae5,
        64'h05130000_3517bae5,
        64'h85930000_359744b0,
        64'h0613a025_04f71e63,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'hb407aa23_00003797,
        64'hc385fd84_3783fcf4,
        64'h262387ba_fcf42823,
        64'h87b2fcf4_2a238736,
        64'h87aefca4_3c230080,
        64'hf822fc06_71398082,
        64'h61457402_70a2853e,
        64'hfec42783_0001fcf7,
        64'h19e301f0_07b7873e,
        64'h27818ff9_01f007b7,
        64'hfe842703_fef42423,
        64'h87aa899f_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'ha839fef4_242387aa,
        64'h8b7fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783fe8f,
        64'he0ef3e80_05139abf,
        64'he0ef853a_02c00593,
        64'h863e93c1_17c20047,
        64'he79393c1_17c2fe44,
        64'h278343d8_fd843783,
        64'hfef42223_87aa999f,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783d3ed,
        64'h27818b89_fe442783,
        64'hfef42223_87aa9b9f,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783a821,
        64'hfef42223_87aa9d1f,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783a1bf,
        64'he0ef853a_02c00593,
        64'h863e93c1_17c20017,
        64'he79393c1_17c2fe44,
        64'h278343d8_fd843783,
        64'hfef42223_87aaa09f,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783a211,
        64'hfef42623_4785e789,
        64'h27818ba1_2781fe24,
        64'h5783fef4_112387aa,
        64'ha33fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'h8c3fe0ef_38878513,
        64'h6785a87f_e0ef853e,
        64'h03e00593_863afe24,
        64'h570343dc_fd843783,
        64'hfef41123_0087e793,
        64'hfe245783_fef41123,
        64'h87aaa75f_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h3783abff_e0ef853e,
        64'h02c00593_863afe24,
        64'h570343dc_fd843783,
        64'hfef41123_9be9fe24,
        64'h5783fef4_112387aa,
        64'haabfe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'hffe12781_8ff901f0,
        64'h07b7fe84_2703fef4,
        64'h242387aa_a33fe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783a839_fef42423,
        64'h87aaa51f_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'hfef42623_4785c781,
        64'h2781fec4_2783fef4,
        64'h262387aa_212000ef,
        64'hfd843503_b0078593,
        64'h67854601_4681fca4,
        64'h3c231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_f3e52781,
        64'h8b892781_feb44783,
        64'hfef405a3_87aabd9f,
        64'he0ef853e_02f00593,
        64'h43dcfd84_3783a821,
        64'hfef405a3_87aabf1f,
        64'he0ef853e_02f00593,
        64'h43dcfd84_3783c3bf,
        64'he0ef853e_02f00593,
        64'h460943dc_fd843783,
        64'hbcdfe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783be3f,
        64'he0ef853a_03000593,
        64'hfff78613_67c143d8,
        64'hfd843783_02e78a23,
        64'h4709fd84_3783a031,
        64'h02e78a23_4705fd84,
        64'h3783c799_2781fec4,
        64'h2783fef4_262387aa,
        64'h2de000ef_fd843503,
        64'h10000593_40ff8637,
        64'h4681a855_fef42623,
        64'h4785a0c1_4785e6e7,
        64'hae234705_00003797,
        64'h99dfe0ef_f0c50513,
        64'h00003517_f0c58593,
        64'h00003597_3ac00613,
        64'ha025cb8d_2781fec4,
        64'h2783fef4_262387aa,
        64'h32e000ef_fd843503,
        64'h45814601_4681ac1f,
        64'he0ef7107_85136789,
        64'hec07a223_00003797,
        64'haa194785_ece7a923,
        64'h47050000_37979f3f,
        64'he0eff625_05130000,
        64'h3517f625_85930000,
        64'h35973ab0_0613a025,
        64'h04f71e63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_f007a423,
        64'h00003797_c385fd84,
        64'h3783fca4_3c231800,
        64'hf022f406_71798082,
        64'h614d64ea_740a70aa,
        64'h853efdc4_27830001,
        64'ha0110001_a0210001,
        64'ha031fcf4_2e234785,
        64'hcb892781_fdc42783,
        64'hfcf42e23_87aa5040,
        64'h10eff584_35032000,
        64'h059302f7_17634785,
        64'h873e0347_c783f584,
        64'h378300f7_1a634791,
        64'h873e57fc_f5843783,
        64'h0001a0b9_fcf42e23,
        64'h4785c791_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h79e020ef_f5843503,
        64'h85befd44_2783fcf4,
        64'h2a231007_879b03a2,
        64'h07b7eb95_0a27c783,
        64'hdb078793_00003797,
        64'ha071fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa09d0,
        64'h10eff584_350302f7,
        64'h11634791_873e57fc,
        64'hf5843783_a865fcf4,
        64'h2e234785_00f70663,
        64'h4785873e_0b97c783,
        64'hdf878793_00003797,
        64'h04f71663_4791873e,
        64'h57fcf584_378300f7,
        64'h09634795_873e57fc,
        64'hf5843783_a8c5fcf4,
        64'h2e234785_00f70663,
        64'h4789873e_0b97c783,
        64'he3078793_00003797,
        64'h02f71063_479d873e,
        64'h57fcf584_3783aa29,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_6ac020ef,
        64'hf5843503_e6458593,
        64'h00003597_a281fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa6570_10eff584,
        64'h35030cf7_0b634799,
        64'h873e57fc_f5843783,
        64'hd7f84719_f5843783,
        64'ha029d7f8_4715f584,
        64'h378300e7_f7634785,
        64'h873e0377_c783f584,
        64'h3783cf91_27818b89,
        64'h27810c47_c783ec67,
        64'h87930000_3797a825,
        64'hd7f84711_f5843783,
        64'h00e7f763_4785873e,
        64'h0377c783_f5843783,
        64'hcf912781_8bb12781,
        64'h0c47c783_ef478793,
        64'h00003797_a09dd7f8,
        64'h471df584_378300e7,
        64'hf7634785_873e0377,
        64'hc783f584_3783cf91,
        64'h27810307_f7932781,
        64'h0c47c783_f2478793,
        64'h00003797_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810d47_c783f3e7,
        64'h87930000_379753f8,
        64'hf5843783_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810087_979b2781,
        64'h0d57c783_f6478793,
        64'h00003797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0107979b_27810d67,
        64'hc783f8a7_87930000,
        64'h379753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b0187_979b2781,
        64'h0d77c783_fac78793,
        64'h00003797_a461fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa01b0_20eff584,
        64'h3503fd25_85930000,
        64'h3597a47d_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h2bf010ef_f5843503,
        64'h28f71263_4795873e,
        64'h0347c783_f5843783,
        64'hacf1fcf4_2e234785,
        64'h28f70d63_4785873e,
        64'h0b97c783_01c78793,
        64'h00003797_ace5fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa08b0_20eff584,
        64'h35030425_85930000,
        64'h3597ae39_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h034020ef_f5843503,
        64'hd7f84715_f5843783,
        64'h2ee7fd63_4785873e,
        64'h0377c783_f5843783,
        64'h30078563_27818b89,
        64'h27810c47_c78308e7,
        64'h87930000_3797d3f8,
        64'hf5843783_0007871b,
        64'h8fd92781_0d47c783,
        64'h0a878793_00003797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h8fd92781_0087979b,
        64'h27810d57_c7830ce7,
        64'h87930000_379753f8,
        64'hf5843783_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810107_979b2781,
        64'h0d67c783_0f478793,
        64'h00003797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_0187979b,
        64'h27810d77_c7831167,
        64'h87930000_3797aecd,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_185020ef,
        64'hf5843503_13c58593,
        64'h00003597_a921fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa4290_10eff584,
        64'h350314f7_1f634785,
        64'h873e0367_c783f584,
        64'h378316e7_f763478d,
        64'h873e0357_c783f584,
        64'h378316f7_1f634789,
        64'h873e0347_c783f584,
        64'h3783a19d_fcf42e23,
        64'h47854207_83632781,
        64'hfdc42783_fcf42e23,
        64'h87aa17e0_20eff584,
        64'h3503d7f8_4715f584,
        64'h378344e7_f3634785,
        64'h873e0377_c783f584,
        64'h37834407_8b632781,
        64'h8b892781_f9d44783,
        64'h46078263_0004c783,
        64'h02e78e23_4705f584,
        64'h3783ff5f_e0ef3e80,
        64'h05139b6f_f0ef853a,
        64'h02c00593_863e93c1,
        64'h17c20047_e793fda4,
        64'h578343d8_f5843783,
        64'hfcf41d23_87aa9a0f,
        64'hf0ef853e_02c00593,
        64'h43dcf584_3783d3e5,
        64'h27818b89_2781fda4,
        64'h5783fcf4_1d2387aa,
        64'h9c2ff0ef_853e02c0,
        64'h059343dc_f5843783,
        64'ha821fcf4_1d2387aa,
        64'h9daff0ef_853e02c0,
        64'h059343dc_f5843783,
        64'ha24ff0ef_853a02c0,
        64'h0593863e_93c117c2,
        64'h0017e793_fda45783,
        64'h43d8f584_3783fcf4,
        64'h1d2387aa_a0eff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_a3a5fcf4,
        64'h2e234785_e7892781,
        64'h8ba12781_fd245783,
        64'hfcf41923_87aaa38f,
        64'hf0ef853e_03e00593,
        64'h43dcf584_37838c8f,
        64'hf0ef3887_85136785,
        64'ha8cff0ef_853e03e0,
        64'h0593863a_fd245703,
        64'h43dcf584_3783fcf4,
        64'h19230087_e793fd24,
        64'h5783fcf4_192387aa,
        64'ha7aff0ef_853e03e0,
        64'h059343dc_f5843783,
        64'hac4ff0ef_853e02c0,
        64'h0593863a_fd245703,
        64'h43dcf584_3783fcf4,
        64'h19239be9_fd245783,
        64'hfcf41923_87aaab0f,
        64'hf0ef853e_02c00593,
        64'h43dcf584_37831407,
        64'h9d6303c7_c783f584,
        64'h378316f7_136347a1,
        64'h873e4bdc_f5843783,
        64'h16e7fa63_478d873e,
        64'hf9d44783_1807d063,
        64'h4187d79b_0187979b,
        64'h0024c783_62079e63,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_18e020ef,
        64'hf5843503_85bef904,
        64'h0793adb9_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h66f010ef_f5843503,
        64'hc3852781_8b912781,
        64'h0014c783_a561fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa4b30_10eff584,
        64'h350385a6_a565fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa34d0_20eff584,
        64'h350326f7_12634785,
        64'h873e0347_c783f584,
        64'h3783add9_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h46c010ef_f5843503,
        64'hadd5fcf4_2e234785,
        64'hadf5fcf4_2e234785,
        64'hcb892781_fdc42783,
        64'hfcf42e23_87aa06f0,
        64'h20eff584_350385be,
        64'h5f9cf584_3783df98,
        64'ha807071b_018cc737,
        64'hf5843783_af05fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa6dc0_10eff584,
        64'h350304f7_1b634795,
        64'h873e0347_c783f584,
        64'h378300f7_0a634789,
        64'h873e0347_c783f584,
        64'h3783a7bd_fcf42e23,
        64'h4785c3d1_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h0e1020ef_f5843503,
        64'h85be5f9c_f5843783,
        64'hdf988407_071b017d,
        64'h8737f584_3783a801,
        64'hdf98ac07_071b0121,
        64'hf737f584_378300f7,
        64'h1a634789_873e0367,
        64'hc783f584_37837c40,
        64'h006ffcf4_2e234785,
        64'hc7912781_fdc42783,
        64'hfcf42e23_87aa915f,
        64'hf0eff584_350306f7,
        64'h1c634785_873e0347,
        64'hc783f584_37837f40,
        64'h006ffcf4_2e234785,
        64'h00f70763_4795873e,
        64'h0347c783_f5843783,
        64'h00f70f63_4789873e,
        64'h0347c783_f5843783,
        64'h02f70763_4785873e,
        64'h0347c783_f5843783,
        64'h02f702e3_47850007,
        64'h871bfdc4_2783fcf4,
        64'h2e2387aa_053000ef,
        64'hf5843503_a83902e7,
        64'h8a234715_f5843783,
        64'h00f71863_400007b7,
        64'h873e2781_8ff9c000,
        64'h07b7873e_579cf584,
        64'h37830750_006f4785,
        64'h7ae7a323_47050000,
        64'h3797ac6f_f0ef8365,
        64'h05130000_45178365,
        64'h85930000_45972400,
        64'h0613a02d_04f71a63,
        64'h4789873e_0367c783,
        64'hf5843783_df98a807,
        64'h071b0006_2737f584,
        64'h37830207_8e23f584,
        64'h378302e7_8a234705,
        64'hf5843783_02e78ba3,
        64'h4705f584_37838007,
        64'ha1230000_47970e10,
        64'h006f4785_80e7a923,
        64'h47050000_4797b32f,
        64'hf0ef8a25_05130000,
        64'h45178a25_85930000,
        64'h459723f0_0613a02d,
        64'h06f71963_11178793,
        64'h111117b7_873e53dc,
        64'hf5843783_8407a423,
        64'h00004797_c385f584,
        64'h3783fc04_3423fc04,
        64'h3023fa04_3c23fa04,
        64'h3823fa04_3423fa04,
        64'h3023f804_3c23f804,
        64'h38230004_b0230057,
        64'h94938395_07fdf807,
        64'h8793fe04_0793f4a4,
        64'h3c231900_ed26f122,
        64'hf5067171_80826161,
        64'h640660a6_853efec4,
        64'h2783fe04_2623d3f8,
        64'hfb843783_0007871b,
        64'h00a7979b_27812785,
        64'h27818ff9_17fd0040,
        64'h07b7873e_27810087,
        64'hd79bfc44_278302f7,
        64'h16634785_873e2781,
        64'h8b8d2781_0167d79b,
        64'hfcc42783_a081d3f8,
        64'hfb843783_0007871b,
        64'h0097d79b_fd042783,
        64'hfcf42823_02f707bb,
        64'hfd842783_fd042703,
        64'hfcf42823_02f707bb,
        64'hfd442703_27812785,
        64'hfd042783_fcf42823,
        64'h8fd9fd04_27830007,
        64'h871b8ff9_c0078793,
        64'h6785873e_278100a7,
        64'h979bfc84_2783fcf4,
        64'h28230167_d79bfc44,
        64'h2783fcf4_2a232781,
        64'h00f717bb_47052781,
        64'h27892781_8b9d2781,
        64'h0077d79b_fc442783,
        64'hfcf42c23_278100f7,
        64'h17bb4705_27818bbd,
        64'h27810087_d79bfc84,
        64'h2783e3c5_27818b8d,
        64'h27810167_d79bfcc4,
        64'h2783fcf4_26232781,
        64'h87aae88f_f0ef853e,
        64'h93811782_278127f1,
        64'h43dcfb84_3783fcf4,
        64'h24232781_87aaea4f,
        64'hf0ef853e_93811782,
        64'h278127e1_43dcfb84,
        64'h3783fcf4_22232781,
        64'h87aaec0f_f0ef853e,
        64'h93811782_278127d1,
        64'h43dcfb84_3783fcf4,
        64'h20232781_87aaedcf,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfb84,
        64'h3783a28d_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h69f000ef_fb843503,
        64'h90078593_6785863e,
        64'h46814bbc_fb843783,
        64'hd7d54bbc_fb843783,
        64'hcbb8fb84_37830007,
        64'h871b8ff9_77c1873e,
        64'h278187aa_f3aff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'ha2c1fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa6fd0,
        64'h00effb84_35033000,
        64'h05934601_4681c7f8,
        64'hfb843783_0007871b,
        64'h87aa81df_f0ef853e,
        64'h45f143dc_fb843783,
        64'hc7b8fb84_37830007,
        64'h871b87aa_837ff0ef,
        64'h853e45e1_43dcfb84,
        64'h3783c3f8_fb843783,
        64'h0007871b_87aa851f,
        64'hf0ef853e_45d143dc,
        64'hfb843783_c3b8fb84,
        64'h37830007_871b87aa,
        64'h86bff0ef_853e45c1,
        64'h43dcfb84_3783a4b9,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_78b000ef,
        64'hfb843503_20000593,
        64'h46014681_ac95fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa5850_00effb84,
        64'h350302e7_8e234705,
        64'hfb843783_c78d2781,
        64'h8ff90100_07b7fe84,
        64'h2703db98_4705fb84,
        64'h3783c789_27818ff9,
        64'h400007b7_fe842703,
        64'hf407dde3_fe842783,
        64'hfef42423_87aa85df,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfb84,
        64'h3783a4cd_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h01e010ef_fb843503,
        64'h90078593_67ad863e,
        64'h4681fe44_2783fef4,
        64'h22238fd9_010007b7,
        64'hfe442703_00f71963,
        64'h47a1873e_4bdcfb84,
        64'h378302f7_10634789,
        64'h873e0367_c783fb84,
        64'h3783fef4_222340ff,
        64'h87b7a689_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h07e010ef_fb843503,
        64'h70078593_678d4601,
        64'h4681a055_fe042423,
        64'h02e78aa3_4709fb84,
        64'h3783a031_02e78aa3,
        64'h4705fb84_378300f7,
        64'h08631aa0_07930007,
        64'h871bfe84_2783fef4,
        64'h242387aa_92bff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'hf3e52781_8b892781,
        64'hfe344783_fef401a3,
        64'h87aaa6df_f0ef853e,
        64'h02f00593_43dcfb84,
        64'h3783a821_fef401a3,
        64'h87aaa85f_f0ef853e,
        64'h02f00593_43dcfb84,
        64'h3783acff_f0ef853e,
        64'h02f00593_460943dc,
        64'hfb843783_04f71863,
        64'h47890007_871bfec4,
        64'h2783a129_fef42623,
        64'h478500f7_06634789,
        64'h0007871b_fec42783,
        64'hcf812781_fec42783,
        64'hfef42623_87aa1540,
        64'h10effb84_35038007,
        64'h85936785_1aa00613,
        64'h4681a189_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h17e010ef_fb843503,
        64'h45814601_4681a19d,
        64'hfef42623_4785e789,
        64'h27818ff9_67c1fdc4,
        64'h2703fcf4_2e2387aa,
        64'ha0fff0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfb84_3783cb8d,
        64'h47dcfb84_378302f7,
        64'h0e634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_fb843783,
        64'ha9754785_d6e7a123,
        64'h47050000_4797883f,
        64'hf0efdf25_05130000,
        64'h4517df25_85930000,
        64'h45971620_0613a025,
        64'h04f71363_4789873e,
        64'h0367c783_fb843783,
        64'hcbd84711_fb843783,
        64'hd807ae23_00004797,
        64'ha3114785_dae7a523,
        64'h47050000_47978cbf,
        64'hf0efe3a5_05130000,
        64'h4517e3a5_85930000,
        64'h45971610_0613a025,
        64'h04f71763_11178793,
        64'h111117b7_873e53dc,
        64'hfb843783_de07a023,
        64'h00004797_c385fb84,
        64'h3783faa4_3c230880,
        64'he0a2e486_715d8082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hbcdff0ef_853e4591,
        64'h20000613_43dcfd84,
        64'h3783e2e7_9223474d,
        64'h00004797_be9ff0ef,
        64'h853e03a0_05934601,
        64'h43dcfd84_3783bfbf,
        64'hf0ef853e_03800593,
        64'h460143dc_fd843783,
        64'hc0dff0ef_853a0360,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c23f,
        64'hf0ef853a_03400593,
        64'heff78613_67c143d8,
        64'hfd843783_cb9ff0ef,
        64'h853e0280_05934661,
        64'h43dcfd84_3783ccbf,
        64'hf0ef853a_02900593,
        64'h863e0ff7_f7930017,
        64'he793feb4_478343d8,
        64'hfd843783_fe0405a3,
        64'ha019fef4_05a347a9,
        64'hc7892781_8ff90400,
        64'h07b7873e_579cfd84,
        64'h3783a005_fef405a3,
        64'h47b1c789_27818ff9,
        64'h020007b7_873e579c,
        64'hfd843783_a82dfef4,
        64'h05a347b9_c7892781,
        64'h8ff90100_07b7873e,
        64'h579cfd84_3783a8d5,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_13c030ef,
        64'hfd843503_a8078593,
        64'h000627b7_b27ff0ef,
        64'h0c800513_00f71663,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cfd84_378302f7,
        64'h13634789_873e0367,
        64'hc783fd84_3783d93f,
        64'hf0ef853e_02900593,
        64'h463d43dc_fd843783,
        64'ha811da7f_f0ef853e,
        64'h02900593_463d43dc,
        64'hfd843783_00f71c63,
        64'h4789873e_0367c783,
        64'hfd843783_d798fd84,
        64'h37830007_871b87aa,
        64'hc7fff0ef_853e9381,
        64'h17822781_0407879b,
        64'h43dcfd84_378302e7,
        64'h8b23fd84_37830ff7,
        64'hf71387aa_d3fff0ef,
        64'h853e0fe0_059343dc,
        64'hfd843783_f3e52781,
        64'h8b852781_fea44783,
        64'hfef40523_87aade1f,
        64'hf0ef853e_02f00593,
        64'h43dcfd84_3783a821,
        64'hfef40523_87aadf9f,
        64'hf0ef853e_02f00593,
        64'h43dcfd84_3783e43f,
        64'hf0ef853e_02f00593,
        64'h460543dc_fd843783,
        64'hc1bff0ef_3e800513,
        64'he5dff0ef_853e0290,
        64'h05934601_43dcfd84,
        64'h3783a811_e71ff0ef,
        64'h853e0290_05934641,
        64'h43dcfd84_3783a481,
        64'h478504e7_a4234705,
        64'h00004797_b69ff0ef,
        64'h0d850513_00004517,
        64'h0d858593_00004597,
        64'h0b500613_a02504f7,
        64'h10634789_873e2781,
        64'h0ff7f793_278187aa,
        64'he03ff0ef_853e0fe0,
        64'h059343dc_fd843783,
        64'h0607b823_fd843783,
        64'hd7f84719_fd843783,
        64'h0607a223_fd843783,
        64'h02e78023_fd843783,
        64'h0207c703_fd043783,
        64'hcfd8fd84_37834fd8,
        64'hfd043783_cf98fd84,
        64'h37834f98_fd043783,
        64'hcbd8fd84_37834bd8,
        64'hfd043783_cb98fd84,
        64'h37834b98_fd043783,
        64'hc7d8fd84_378347d8,
        64'hfd043783_d3d81117,
        64'h071b1111_1737fd84,
        64'h3783c798_fd843783,
        64'h4798fd04_3783c3d8,
        64'hfcc42703_fd843783,
        64'h00e79023_fd843783,
        64'h0007d703_fd043783,
        64'h1207a223_00004797,
        64'ha62d4785_12e7a923,
        64'h47050000_4797c53f,
        64'hf0ef1c25_05130000,
        64'h45171c25_85930000,
        64'h45970b40_0613a025,
        64'hc7fdfd04_37831407,
        64'had230000_4797cb89,
        64'hfd843783_fcf42623,
        64'h87b2fcb4_3823fca4,
        64'h3c230080_f822fc06,
        64'h71398082_61056442,
        64'h60e20001_e8dff0ef,
        64'h853e85ba_fea44703,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_052387ba,
        64'hfef405a3_87b6fef4,
        64'h26238732_86ae87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h853e87aa_e7fff0ef,
        64'h853e9381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef405a3,
        64'h87bafef4_2623872e,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e20001_f39ff0ef,
        64'h853e85ba_fe845703,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_142387ba,
        64'hfef405a3_87b6fef4,
        64'h26238732_86ae87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h853e87aa_f1dff0ef,
        64'h853e9381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef405a3,
        64'h87bafef4_2623872e,
        64'h87aa1000_e822ec06,
        64'h11018082_61457422,
        64'h0001c398_fd442703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf42a23,
        64'h87aefca4_3c231800,
        64'hf4227179_80826145,
        64'h74220001_00e79023,
        64'hfd645703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf41b23_87aefca4,
        64'h3c231800_f4227179,
        64'h80826145_74220001,
        64'h00e78023_fd744703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf40ba3,
        64'h87aefca4_3c231800,
        64'hf4227179_80826105,
        64'h6462853e_2781439c,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61056462_853e93c1,
        64'h17c20007_d783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826105,
        64'h6462853e_0ff7f793,
        64'h0007c783_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61457422,
        64'h853efe84_3783fae7,
        64'hf5e34785_0007871b,
        64'hfe442783_fef42223,
        64'h2785fe44_2783a829,
        64'hfef43423_97baefe7,
        64'h07130000_4717078a,
        64'h97ba078e_87bafe44,
        64'h670302f7_10632781,
        64'h2701fde4_57030007,
        64'hd78397ba_f3068713,
        64'h078a97ba_078e87ba,
        64'hfe446703_00004697,
        64'ha0b9fe04_2223fe04,
        64'h3423fcf4_1f2387aa,
        64'h1800f422_71798082,
        64'hfea7ede3_8f99ff86,
        64'hb7830200_c6b702f5,
        64'h05330280_0793fee7,
        64'h8ee3ff86_b7030200,
        64'hc6b7ff87_b7830200,
        64'hc7b78082_ff87b503,
        64'h0200c7b7_80826125,
        64'h70a2a1bf_f0efe43a,
        64'hecc6e8c2_e4bef406,
        64'h72c50513_567d080c,
        64'h86b21838_ec2ee0ba,
        64'hfc36ffff_f517e82a,
        64'h711da43f_f06f72e5,
        64'h0513ffff_f51785aa,
        64'h862e86b2_87368082,
        64'h610560e2_a5dff0ef,
        64'hec06a645_0513002c,
        64'h567d872e_00000517,
        64'h86aa1101_80826161,
        64'h60e2a7bf_f0efe43a,
        64'he4c6e0c2_fc3eec06,
        64'h10387745_0513f83a,
        64'hfffff517_85aa862e,
        64'h86b2f436_715d8082,
        64'h616160e2_aa5ff0ef,
        64'he43ae4c6_e0c2fc3e,
        64'hec067a25_05131018,
        64'h567df83a_f032ffff,
        64'hf51785aa_86aef436,
        64'h715d8082_612560e2,
        64'had1ff0ef_e43aecc6,
        64'he8c2e4be_ec06ae65,
        64'h0513567d_1038858a,
        64'he0baf832_f42e0000,
        64'h051786aa_fc36711d,
        64'hb31d4809_b32d4821,
        64'hbb1d4841_0206e693,
        64'hbb498da2_99020250,
        64'h051385d2_866e86ce,
        64'h001d8413_b7d58622,
        64'h2c859902_00160413,
        64'h02000513_85d286ce,
        64'hbb6d8db2_8aea018c,
        64'he563c019_fc089de3,
        64'hfff8869b_fe0a82e3,
        64'hc51901b7_06330007,
        64'h450378a2_77029902,
        64'h85d286ce_f83af03a,
        64'hf4460705_88b6b7e1,
        64'h78c28df2_8cc27762,
        64'h7e027822_99020200,
        64'h051385d2_86ce866e,
        64'hf072f442_f846fc3a,
        64'h001d8e13_b7c90785,
        64'ha08140ed_8db38cc2,
        64'h018ce863_001c881b,
        64'he4110006_841b8a89,
        64'h00060c9b_8666011c,
        64'hf3638646_000a8863,
        64'h40e78cbb_2a814006,
        64'hfa9302f6_1b63c199,
        64'h0007c583_87ba00f7,
        64'h06339381_02089793,
        64'h00088563_57fd000a,
        64'hb703008a_8d13b7cd,
        64'h8ca22b05_99020200,
        64'h051385d2_86ce001c,
        64'h84138666_b5598de6,
        64'h8aea018b_6563c019,
        64'h9902001d_8c93008a,
        64'h8d1385d2_866e86ce,
        64'h000ac503_ff8764e3,
        64'h001d8d13_00170b1b,
        64'h8dea875a_99020200,
        64'h051385d2_86ce866e,
        64'ha8094705_e00d4b05,
        64'h0006841b_8a89b7ed,
        64'h8f7d67e2_dbe50807,
        64'hf793b769_93014781,
        64'he062e436_17020ff7,
        64'h7713ca09_000aa703,
        64'h0407f613_b755e062,
        64'he4364781_000ab703,
        64'hc7191007_f713bde5,
        64'h4781e062_e436000a,
        64'hb703c719_bff1000a,
        64'ha783b7cd_000a9783,
        64'hc7810807_f793bfd9,
        64'h40e6073b_93fde062,
        64'he43600e7_c63341f7,
        64'hd71b000a_c783cf09,
        64'h0406f713_b789bb7f,
        64'hf0ef854a_85d2866e,
        64'h86ce93fd_40e60733,
        64'h00f74633_43f7d713,
        64'he062e436_000ab783,
        64'hc31d87b6_1006f713,
        64'hb5dd0780_0793eef5,
        64'h09e30750_0793a89d,
        64'h4841e03e_e436008a,
        64'h8413000a_b70347c1,
        64'h0216e693_d4f51ae3,
        64'h07000793_f0f50ce3,
        64'h06f00793_02a7e563,
        64'h12f50f63_07300793,
        64'hb71d0640_07930ef5,
        64'h06630630_0793bddd,
        64'h0c06e693_8082614d,
        64'h6da66d46_6ce67c06,
        64'h7ba67b46_7ae66a0a,
        64'h69aa694a_64ea000d,
        64'h851b740a_70aa9902,
        64'h450185d2_86cefff9,
        64'h8613013d_e463866e,
        64'hda0517e3_0004c503,
        64'h8aa28daa_cf5ff0ef,
        64'h854a85d2_866e86ce,
        64'h93fd40e6_073300f7,
        64'h463343f7_d713e062,
        64'he436000a_b783cf45,
        64'h10c51c63_06400613,
        64'h00c50663_008a8413,
        64'h02085813_270187b6,
        64'h06900613_18022006,
        64'hf7139af9_c3914006,
        64'hf7939acd_00f50363,
        64'h06400793_00f50763,
        64'h48299abd_06900793,
        64'h2ef50463_06200793,
        64'h2ef50663_06f00793,
        64'h2ef50663_05800793,
        64'h2ef50c63_07800793,
        64'he4f514e3_05800793,
        64'h2ef50863_02500793,
        64'h0ca7ef63_00f50c63,
        64'h06200793_0ea7ec63,
        64'h02f50263_00170493,
        64'h06900793_00074503,
        64'h0806e693_0ef60e63,
        64'h0014c603_a0390024,
        64'h87133006_e693a821,
        64'h1006e693_00f60563,
        64'h0014c603_b7e907a0,
        64'h061300c7_89630740,
        64'h0613bf65_84babf75,
        64'h8abe0489_28814881,
        64'h0008d363_008a8793,
        64'h000aa883_00f61d63,
        64'h02a00793_a8998726,
        64'h04c78063_06a00613,
        64'h04c78c63_06800613,
        64'h02f66d63_04c78663,
        64'h00148713_06c00613,
        64'h0004c783_fef671e3,
        64'h0ff7f793_fd07079b,
        64'h00148593_0004c703,
        64'h00e888bb_fd08889b,
        64'h84ae031b_88bbb775,
        64'h84b28aba_40f00c3b,
        64'h0026e693_0007d663,
        64'h00078c1b_008a8713,
        64'h000aa783_fce796e3,
        64'h4c0102a0_0713a825,
        64'h462584ba_06f5ee63,
        64'h4006e693_0ff7f793,
        64'hfd06079b_00148713,
        64'h45a50014_c60306f7,
        64'h17634881_02e00793,
        64'h0004c703_fef671e3,
        64'h0ff7f793_fd07079b,
        64'h00148593_0004c703,
        64'h00e30c3b_fd03031b,
        64'h84ae038b_833bbf75,
        64'h0106e693_b7c90086,
        64'he693b7e1_0046e693,
        64'hb7f90026_e693a025,
        64'h46254c01_06e5e963,
        64'h45a50ff7_7713fd07,
        64'h871b02a7_856302b7,
        64'h8463fcf7_6fe302e7,
        64'h85630014_86130004,
        64'hc78384b2_0016e693,
        64'h02879163_03000413,
        64'h02878f63_02d00413,
        64'ha8210230_05130200,
        64'h059302b0_07134681,
        64'ha15585d2_866e86ce,
        64'h001d8413_00f50863,
        64'h04850250_0793ac81,
        64'h4ba9ec3e_4d81fffb,
        64'h07936b41_cc890913,
        64'h00000917_e589892a,
        64'h8aba84b6_89b28a2e,
        64'he4eee8ea_ece6f0e2,
        64'hf4def8da_f122f506,
        64'hfcd6e152_e54ee94a,
        64'hed267171_808298df,
        64'hf06fc119_b7e1006e,
        64'h033b8082_616160a6,
        64'hd17ff0ef_887e1018,
        64'h0008089b_e43ae876,
        64'he0464746_fc579de3,
        64'hc319fe6f_0fa39f3e,
        64'h0ff37313_02010f13,
        64'h07850307_57330303,
        64'h031b03e3_ee630fff,
        64'h73130307_7f330200,
        64'h0293ff63_0e1b43a5,
        64'h47810410_0313000e,
        64'h04630610_0313020e,
        64'hfe13c721_47810003,
        64'h0463400e_f313fefe,
        64'hfe93e319_4ee68fbe,
        64'he486715d_b7e1006e,
        64'h033b8082_616160a6,
        64'hd97ff0ef_887e1018,
        64'h0008089b_e43ae876,
        64'he0464746_fc579de3,
        64'hc319fe6f_0fa39f3e,
        64'h0ff37313_02010f13,
        64'h07850307_57330303,
        64'h031b03e3_ee630fff,
        64'h73130307_7f330200,
        64'h0293ff63_0e1b43a5,
        64'h47810410_0313000e,
        64'h04630610_0313020e,
        64'hfe13c721_47810003,
        64'h0463400e_f313fefe,
        64'hfe93e319_4ee68fbe,
        64'he486715d_b7a98622,
        64'h9b020016_04130200,
        64'h051385de_86e2b791,
        64'h9b0285de_86e20009,
        64'h4503b7ed_41540cb3,
        64'h02095913_02099913,
        64'hbf89ff27_e3e3009c,
        64'h87b384ea_00148d13,
        64'h67229b02_e43a0200,
        64'h051385de_86e28626,
        64'hb7ad00d6_00230087,
        64'h0633da3d_0087f613,
        64'hbf9d02b0_06130087,
        64'h06b3c611_0047f613,
        64'hbfa10620_06130087,
        64'h06b3f886_ece346fd,
        64'hf6d898e3_4689b7bd,
        64'h05800613_008706b3,
        64'hfa86e7e3_46fd8082,
        64'h61658532_6d426ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_0b37e163,
        64'h415607b3_0209d993,
        64'h1982000a_09630094,
        64'h06330b2c_9663197d,
        64'h412d0633_01248d33,
        64'hfff70c93_00870933,
        64'hcbcd84d6_8b8d0405,
        64'h00c68023_02d00613,
        64'h008706b3_08080463,
        64'h00d40b63_02000693,
        64'h040500c6_80230300,
        64'h06130087_06b30286,
        64'he66346fd_040500c6,
        64'h80230780_06130087,
        64'h06b30486_e06346fd,
        64'head10207_f6930ad8,
        64'h966346c1_4401bf55,
        64'hfe6e0fa3_00870e33,
        64'h0405a0e9_02c89a63,
        64'h84364609_02c88163,
        64'h14794641_c285fff4,
        64'h06930286_95639281,
        64'h02099693_00868763,
        64'h92811682_cc0dee15,
        64'h4007f613_ca3d0107,
        64'hf61302b4_1e6300a4,
        64'h7463c609_03000313,
        64'h02000593_91010209,
        64'h9513fea4_69e3fe6e,
        64'h0fa30087_0e330405,
        64'h00b40963_a8010300,
        64'h03130200_05939101,
        64'h02069513_39fdc191,
        64'h00c7f593_00081563,
        64'hc6190009_89630017,
        64'hf613040a_1a6359e6,
        64'h56c68ab2_8bae8b2a,
        64'h8c362a01_e86aec66,
        64'he8caeca6_f486f062,
        64'hf45ef85a_fc560027,
        64'hfa13e4ce_e0d2478a,
        64'h843ef0a2_71598082,
        64'h8302658c_0005b303,
        64'hc5098082_808200a5,
        64'h802395b2_00d67563,
        64'hbbe102f0_00efd7e5,
        64'h05130000_6517bd35,
        64'hb4250513_85a60000,
        64'h65170470_00efb365,
        64'h05130000_6517cd09,
        64'h84aada9f_f0ef8552,
        64'h865a020a_a5830630,
        64'h00efd9a5_05130000,
        64'h6517f579_90e30804,
        64'h84930770_00ef2985,
        64'ha8850513_00006517,
        64'hff2c17e3_089000ef,
        64'h0905d3a5_05130000,
        64'h65170009_45830704,
        64'h8c130284_89130a30,
        64'h00efdc25_05130000,
        64'h65170af0_00efdb65,
        64'h05130000_6517708c,
        64'h0bd000ef_dac50513,
        64'h00006517_6c8c0cb0,
        64'h00efda25_05130000,
        64'h6517688c_ff2c17e3,
        64'h0dd000ef_0905d8e5,
        64'h05130000_65170009,
        64'h45830109_0c130f30,
        64'h00efdaa5_05130000,
        64'h6517fe99_17e31030,
        64'h00ef0905_db450513,
        64'h00006517_00094583,
        64'hff048913_119000ef,
        64'hda850513_00006517,
        64'h125000ef_d9e50513,
        64'h85ce0000_6517bf15,
        64'hd8a50513_85ce0000,
        64'h651713f0_00efc2e5,
        64'h05130000_6517cd09,
        64'h4b910804_89aa8a8a,
        64'hea7ff0ef_850a4605,
        64'h710144ac_161000ef,
        64'hd9850513_00006517,
        64'h45d616f0_00efd865,
        64'h05130000_651745c6,
        64'h17d000ef_d6c50513,
        64'h00006517_65a618b0,
        64'h00efd625_05130000,
        64'h65177582_199000ef,
        64'hd5850513_00006517,
        64'h65e21a70_00efd4e5,
        64'h05130000_651745d2,
        64'h1b5000ef_d4450513,
        64'h00006517_45c21c30,
        64'h00efd3a5_05130000,
        64'h651745b2_1d1000ef,
        64'hd3050513_00006517,
        64'h45a21df0_00efd265,
        64'h05130000_65176582,
        64'h1ed000ef_d1450513,
        64'h00006517_b75554f9,
        64'h1fd000ef_d0450513,
        64'h00006517_fa843583,
        64'h20d000ef_cfc50513,
        64'h00006517_faa43423,
        64'hc11df71f_f0ef848a,
        64'h850a4585_46057101,
        64'h22d000ef_d0450513,
        64'h00006517_80826125,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h64468526_60e6fa04,
        64'h011354fd_259000ef,
        64'hd0850513_00006517,
        64'hc51df39f_f0ef8b2e,
        64'h8a2a1080_e862ec5e,
        64'hf456fc4e_e0cae4a6,
        64'hec86f05a_f852e8a2,
        64'h711d8082_014160a2,
        64'h557d28f0_00efd1e5,
        64'h05130000_651785aa,
        64'hc90922b0_20efe406,
        64'hc0c50513_46051141,
        64'h00005517_86aab76d,
        64'h45012b70_00efd265,
        64'h05130000_6517bf6d,
        64'h55752c70_00efd065,
        64'h05130000_6517c909,
        64'h85aa1c80_10ef8522,
        64'hbfd15579_2e1000ef,
        64'hcf850513_00006517,
        64'hc90985aa_65f000ef,
        64'h852285aa_c5c40413,
        64'h00005417_41508082,
        64'h01416402_60a2557d,
        64'h30d000ef_d0450513,
        64'h00006517_ed014350,
        64'h00ef4501_321000ef,
        64'he022e406_d0650513,
        64'h11410000_65178082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_00a78223,
        64'h0ff57513_00d78023,
        64'h0085551b_0ff57693,
        64'h00d78623_f8000693,
        64'h00078223_01e71793,
        64'h470d02b5_553b0045,
        64'h959b8082_00a78023,
        64'hdf650207_77130147,
        64'hc70307fa_478d8082,
        64'h02057513_0147c503,
        64'h07fa478d_80820005,
        64'h45038082_00b50023,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_100004b7,
        64'h1c858593_00005597,
        64'hf1402573_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_423040ef,
        64'h40000137_03249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
