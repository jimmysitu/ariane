/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 3895;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_20000060,
        64'h00000000_20000060,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0000000b_0005deec,
        64'he66d1234_abcd330e,
        64'h00000000_00000001,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_200006f8,
        64'h00000000_20000648,
        64'h00000000_20000598,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000030_00003000,
        64'h00000020_00002000,
        64'h00000010_00001000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_322d746c,
        64'h75616665_642d6972,
        64'h742c786e_6c780074,
        64'h6c756166_65642d69,
        64'h72742c78_6e6c7800,
        64'h6c617564_2d73692c,
        64'h786e6c78_00746e65,
        64'h73657270_2d747075,
        64'h72726574_6e692c78,
        64'h6e6c7800_68746469,
        64'h772d326f_6970672c,
        64'h786e6c78_00687464,
        64'h69772d6f_6970672c,
        64'h786e6c78_00322d74,
        64'h6c756166_65642d74,
        64'h756f642c_786e6c78,
        64'h00746c75_61666564,
        64'h2d74756f_642c786e,
        64'h6c780032_2d737475,
        64'h706e692d_6c6c612c,
        64'h786e6c78_00737475,
        64'h706e692d_6c6c612c,
        64'h786e6c78_0072656c,
        64'h6c6f7274_6e6f632d,
        64'h6f697067_00736c6c,
        64'h65632d6f_69706723,
        64'h0070772d_656c6261,
        64'h73696400_7365676e,
        64'h61722d65_6761746c,
        64'h6f760079_636e6575,
        64'h71657266_2d78616d,
        64'h2d697073_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_5a020000,
        64'h04000000_03000000,
        64'hffffffff_49020000,
        64'h04000000_03000000,
        64'h01000000_3c020000,
        64'h04000000_03000000,
        64'h00000000_25020000,
        64'h04000000_03000000,
        64'h08000000_14020000,
        64'h04000000_03000000,
        64'h08000000_04020000,
        64'h04000000_03000000,
        64'h00000000_f0010000,
        64'h04000000_03000000,
        64'h00000000_de010000,
        64'h04000000_03000000,
        64'h00000000_cc010000,
        64'h04000000_03000000,
        64'h00000000_bc010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h000000c1_00000000,
        64'h67000000_10000000,
        64'h03000000_ac010000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'ha0010000_04000000,
        64'h03000000_00000030,
        64'h30303030_30316340,
        64'h6f697067_01000000,
        64'h02000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_03000000,
        64'h52010000_04000000,
        64'h03000000_00000000,
        64'h64656c62_61736964,
        64'h6b000000_09000000,
        64'h03000000_00100000,
        64'h00000000_00b000e0,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00006d65_672c736e,
        64'h6463006d_65672d71,
        64'h6e797a2c_736e6463,
        64'h1b000000_17000000,
        64'h03000000_00000030,
        64'h30306230_30306540,
        64'h74656e72_65687465,
        64'h01000000_02000000,
        64'h02000000_95010000,
        64'h00000000_03000000,
        64'he40c0000_e40c0000,
        64'h86010000_08000000,
        64'h03000000_20bcbe00,
        64'h74010000_04000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00000000,
        64'h746f6c73_2d697073,
        64'h2d636d6d_1b000000,
        64'h0d000000_03000000,
        64'h00000030_40636d6d,
        64'h01000000_00100000,
        64'h00000000_000010e0,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_52010000,
        64'h04000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h00000000_64656c62,
        64'h61736964_6b000000,
        64'h09000000_03000000,
        64'h00000061_392e382d,
        64'h69636864_732c6e61,
        64'h73617261_1b000000,
        64'h12000000_03000000,
        64'h00000000_30303030,
        64'h30313065_40636d6d,
        64'h01000000_02000000,
        64'h00100000_00000000,
        64'h00d000e0_00000000,
        64'h67000000_10000000,
        64'h03000000_02000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h64656c62_61736964,
        64'h6b000000_09000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_0000302e,
        64'h312d6970_73712d71,
        64'h6e797a2c_786e6c78,
        64'h1b000000_13000000,
        64'h03000000_00000000,
        64'h30303064_30303065,
        64'h40697073_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_005a6202,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_000000c0,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30306340,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000030_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h31407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_005a6202,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30634074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08090000_6d020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h40090000_38000000,
        64'had0b0000_edfe0dd0,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'hffffb124_ffffb7c0,
        64'hffffb7c0_ffffb124,
        64'hffffb7c0_ffffb5aa,
        64'hffffb7c0_ffffb7c0,
        64'hffffb6e4_ffffb124,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb124,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb124_ffffb4e6,
        64'hffffb124_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb124_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb7c0,
        64'hffffb7c0_ffffb794,
        64'hffffb10e_ffffb126,
        64'hffffb126_ffffb126,
        64'hffffb126_ffffb126,
        64'hffffb0de_ffffb126,
        64'hffffb126_ffffb126,
        64'hffffb126_ffffb126,
        64'hffffb126_ffffb126,
        64'hffffb05e_ffffb126,
        64'hffffb0f6_ffffb126,
        64'hffffb09e_ffffaeaa,
        64'hffffaf40_ffffaf40,
        64'hffffaec8_ffffaf40,
        64'hffffaee6_ffffaf40,
        64'hffffaf40_ffffaf40,
        64'hffffaf40_ffffaf40,
        64'hffffaf40_ffffaf40,
        64'hffffaf22_ffffaf40,
        64'hffffaf40_ffffaf04,
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00586c6c_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000000_00007525,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000000_00007525,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_58323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h000a5838_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h000a5838_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_000a586c,
        64'h6c363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h00000000_0a756c6c,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h00000000_0a756c6c,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_0a583830,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_0a583830,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_0a583830,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_0a583830,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h00000000_0000000a,
        64'h00000000_00006325,
        64'h00202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h00000000_0a642520,
        64'h3a737574_61747320,
        64'h2c64656c_69616620,
        64'h64616552_20304453,
        64'h00000000_0a216465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a6425,
        64'h203a7375_74617473,
        64'h202c6465_6c696166,
        64'h206e6f69_74617a69,
        64'h6c616974_696e6920,
        64'h64726163_20304453,
        64'h0000000a_6425203a,
        64'h73757461_7473202c,
        64'h64656c69_6166206c,
        64'h61697469_6e692067,
        64'h69666e6f_63204453,
        64'h00000000_0000000a,
        64'h2164656c_69616620,
        64'h6769666e_6f632070,
        64'h756b6f6f_6c204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000020_58323025,
        64'h00000000_0000000a,
        64'h786c6c25_78304045,
        64'h5341425f_4d415244,
        64'h00000000_0000000a,
        64'h000a6425_202c6425,
        64'h00000000_002e2e2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00010198,
        64'h00000000_000101d8,
        64'h00000000_80827b07,
        64'hb5032000_07b7a001,
        64'ha001c100_00a000ef,
        64'h4080043b_e406842a,
        64'he0221141_00055c63,
        64'h00000073_05d00893,
        64'h47814701_46814601,
        64'h4581bfc9_9682852e,
        64'hbfe19682_8556e781,
        64'h27818ff1_11093583,
        64'h31442783_bfd90009,
        64'h3823bf49_fcf406e3,
        64'hf9771de3_1f89b783,
        64'h44189682_ef092701,
        64'h8f710084_2b83009b,
        64'h163b3104_2703d6f5,
        64'hc4040297_966337fd,
        64'h01093683_441cbfd9,
        64'h196134fd_01478563,
        64'h21093783_000a0963,
        64'h80826161_6ba26b42,
        64'h6ae27a02_79a27942,
        64'h74e26406_60a60004,
        64'hdd639922_00349913,
        64'h34fd4404_c8011f89,
        64'hb4034b05_8a2e8aaa,
        64'he45ef84a_fc26e0a2,
        64'he486e85a_ec56f052,
        64'h7a87b983_f44e2000,
        64'h07b7715d_80824501,
        64'he38c97ba_c794070e,
        64'h07090017_069b30c7,
        64'haa238e55_3147a683,
        64'h00d31763_468920d8,
        64'h38233117_a82300c8,
        64'he8b300e6_163b4605,
        64'h3107a883_10c83823,
        64'h983e0037_18130203,
        64'h0a6304e8_4463557d,
        64'h487d4798_1ef73c23,
        64'h20070793_e7891f87,
        64'h3783832a_7a87b703,
        64'h200007b7_b79df8c3,
        64'h71e3963e_8f1d17c1,
        64'h8096fa26_80e78286,
        64'h96960000_02970027,
        64'h9693b759_8dd50205,
        64'h96938dd5_01059693,
        64'h8dd50085_96930ff5,
        64'hf5938082_00b70023,
        64'h00b700a3_00b70123,
        64'h00b701a3_00b70223,
        64'h00b702a3_00b70323,
        64'h00b703a3_00b70423,
        64'h00b704a3_00b70523,
        64'h00b705a3_00b70623,
        64'h00b706a3_00b70723,
        64'h00a68067_96960000,
        64'h0297068a_40c306b3,
        64'h8082e211_fed76de3,
        64'h0741e70c_e30c96ba,
        64'h8a3dff06_7693e1bd,
        64'he3c100f7_779302c3,
        64'h7163872a_433dbff9,
        64'h978204a1_0905609c,
        64'hb7e99782_04a10905,
        64'h609c8082_61056902,
        64'h64a26442_60e20089,
        64'h1d634901_fb848493,
        64'h840d8c1d_fc040413,
        64'hfb848793_6459bc0f,
        64'ha0ef64d9_02891763,
        64'h4901fb44_8493840d,
        64'hec06e04a_8c1dfb44,
        64'h0413fb44_879364d9,
        64'h6459e426_e8221101,
        64'hbff99782_ff87b783,
        64'h97ca0485_033487b3,
        64'hbfafa06f_614569a2,
        64'h694264e2_70a27402,
        64'h00941a63_59e1fc87,
        64'h89134481_840df406,
        64'he44ee84a_ec268c19,
        64'hfc878413_fc070713,
        64'hf0226759_67d97179,
        64'h272000ef_85229782,
        64'hc3916d3c_7a87b503,
        64'h200007b7_1d4000ef,
        64'h842ae406_e0224581,
        64'h114117a0_006f4501,
        64'h46014681_85aa8082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'ha14fc0ef_4505a031,
        64'hfef42623_4785e789,
        64'h27810807_f7932781,
        64'h87aaaa5f_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h37830001_a011f6e7,
        64'hfee30270_07930ff7,
        64'hf713fe94_4783fef4,
        64'h04a32785_fe944783,
        64'hcf992781_0407f793,
        64'h278187aa_adffe0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_a0adfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaae5f_d0effd84,
        64'h35035007_85936785,
        64'h46014685_a829fef4,
        64'h262387aa_afffd0ef,
        64'hfd843503_30078593,
        64'h67854601_468500f7,
        64'h1f634785_873e0347,
        64'hc783fd84_3783a8ad,
        64'hfe0404a3_ad0fc0ef,
        64'h4505b87f_e0ef853e,
        64'h03e00593_863afe64,
        64'h570343dc_fd843783,
        64'hfef41323_0407e793,
        64'hfe645783_fef41323,
        64'h87aab75f_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h3783c2e1_90234741,
        64'hbc5fe0ef_853e4591,
        64'h863afea4_570343dc,
        64'hfd843783_fef41523,
        64'h8ff917fd_6785fea4,
        64'h5703fef4_15230017,
        64'h979bfea4_5783aa25,
        64'h4785c0e1_ae234705,
        64'h93afc0ef_a8450513,
        64'h00001517_a7c58593,
        64'h00001597_4b600613,
        64'ha01502f7_1a63478d,
        64'h873e0377_c783fd84,
        64'h3783fef4_15230400,
        64'h0793c001_ae23aaa5,
        64'h4785c0e1_ae234705,
        64'h97afc0ef_ac450513,
        64'h00001517_abc58593,
        64'h00001597_4b500613,
        64'ha01504f7_13631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783c001,
        64'hae23cf91_fd843783,
        64'hfca43c23_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aabeff,
        64'he0ef853e_93811782,
        64'h278127c1_43dcfd84,
        64'h3783caff_e0ef853e,
        64'h03000593_460943dc,
        64'hfd843783_dfc52781,
        64'h8b89fe84_2783a83d,
        64'hfef42623_4785cd3f,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c3852781,
        64'h8ff967a1_fe842703,
        64'hfef42423_87aacc1f,
        64'he0ef853e_03000593,
        64'h43dcfd84_3783a8bd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_cc7fd0ef,
        64'hfd843503_60000593,
        64'h863e4681_fd442783,
        64'hfcf42a23_87aefca4,
        64'h3c231800_f022f406,
        64'h71798082_61217442,
        64'h70e2853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_cb5fe0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fc843783,
        64'hd75fe0ef_853e0300,
        64'h05934609_43dcfc84,
        64'h3783dfc5_27818b89,
        64'hfdc42783_a83dfef4,
        64'h26234785_d99fe0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fc84,
        64'h3783c385_27818ff9,
        64'h67a1fdc4_2703fcf4,
        64'h2e2387aa_d87fe0ef,
        64'h853e0300_059343dc,
        64'hfc843783_a8bdfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aad8df_d0effc84,
        64'h35038007_85936785,
        64'h863e4685_fe442783,
        64'hc2e19023_47457010,
        64'hd0737010_50730ff0,
        64'h000ffc2f_e0effc84,
        64'h350385be_fc043603,
        64'h2781fe24_5783e23f,
        64'he0ef853e_4591863a,
        64'hfe045703_43dcfc84,
        64'h3783fef4_10238ff9,
        64'h17fd6785_fe045703,
        64'hfef41023_20000793,
        64'hfef41123_4785fce7,
        64'hdee31ff0_07930007,
        64'h871bfe84_2783fef4,
        64'h24232785_fe842783,
        64'h00078023_97bafc04,
        64'h3703fe84_2783a235,
        64'h4785c0e1_ae234705,
        64'hbc2fc0ef_d0c50513,
        64'h00001517_d0458593,
        64'h00001597_37500613,
        64'ha835fe04_2423c001,
        64'hae23aaa1_4785c0e1,
        64'hae234705_beefc0ef,
        64'hd3850513_00001517,
        64'hd3058593_00001597,
        64'h37400613_a01502f7,
        64'h19631117_87931111,
        64'h17b7873e_53dcfc84,
        64'h3783c001_ae23cf91,
        64'hfc843783_fe042223,
        64'hfcb43023_fca43423,
        64'h0080f822_fc067139,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623a019_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hecbfd0ef_fd843503,
        64'ha0078593_67ad4601,
        64'h4681a03d_fef42623,
        64'h4785a82d_4785c0e1,
        64'hae234705_c86fc0ef,
        64'hdd050513_00001517,
        64'hdc858593_00001597,
        64'h34500613_a015c79d,
        64'h2781fec4_2783fef4,
        64'h262387aa_f17fd0ef,
        64'hfd843503_70078593,
        64'h678d863e_46814bbc,
        64'hfd843783_c001ae23,
        64'ha0614785_c0e1ae23,
        64'h4705cd4f_c0efe1e5,
        64'h05130000_1517e165,
        64'h85930000_15973440,
        64'h0613a015_04f71a63,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'hc001ae23_cf91fd84,
        64'h3783fca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'hfe842783_fe042423,
        64'hfedfe0ef_853a02c0,
        64'h0593863e_93c117c2,
        64'h0047e793_fe445783,
        64'h43d8fd84_3783fef4,
        64'h122387aa_fd7fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_d3e52781,
        64'h8b892781_fe645783,
        64'hfef41323_87aaff9f,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783a821,
        64'hfef41323_87aa810f,
        64'hf0ef853e_02c00593,
        64'h43dcfd84_378385af,
        64'hf0ef853e_02c00593,
        64'h863afe44_570343dc,
        64'hfd843783_fef41223,
        64'h0017e793_93c117c2,
        64'h8fd9fe44_5783fec4,
        64'h5703fef4_1623f007,
        64'hf793fec4_5783fef4,
        64'h16230087_979bfec4,
        64'h5783fef4_12230ff7,
        64'hf793fe44_5783fef4,
        64'h122387aa_876ff0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a0a58c2f,
        64'hf0ef853e_02c00593,
        64'h863afe44_570343dc,
        64'hfd843783_fef41223,
        64'h0017e793_93c117c2,
        64'h8fd9fe44_57839341,
        64'h03079713_8fd9fe24,
        64'h5783fec4_5703fef4,
        64'h1623f007_f793fec4,
        64'h5783fef4_16230087,
        64'h979bfec4_5783fef4,
        64'h11230c07_f793fe24,
        64'h5783fef4_11230067,
        64'h979bfe24_5783fef4,
        64'h11230087_d79bfec4,
        64'h5783fef4_122303f7,
        64'hf793fe44_5783fef4,
        64'h122387aa_90eff0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_08f71e63,
        64'h4789873e_0367c783,
        64'hfd843783_a249fef4,
        64'h24234785_00e7f663,
        64'h10000793_0007871b,
        64'hfee45783_fae7fee3,
        64'h10000793_0007871b,
        64'hfee45783_fef41723,
        64'h0017979b_fee45783,
        64'ha839fef4_16230017,
        64'hd79bfee4_578300e7,
        64'he9632781_fd442783,
        64'h0007871b_02f757bb,
        64'h2781fee4_57834798,
        64'hfd843783_a82dfef4,
        64'h17234785_a2edfef4,
        64'h24234785_06e7fa63,
        64'h7fe00793_0007871b,
        64'hfee45783_fae7ffe3,
        64'h7fe00793_0007871b,
        64'hfee45783_fef41723,
        64'h2785fee4_5783a831,
        64'hfef41623_0017d79b,
        64'hfee45783_00e7e963,
        64'h2781fd44_27830007,
        64'h871b02f7_57bb2781,
        64'hfee45783_4798fd84,
        64'h3783a825_fef41723,
        64'h4785ac91_4785c0e1,
        64'hae234705_f7efc0ef,
        64'h0c850513_00001517,
        64'h0c058593_00001597,
        64'h2d000613_a01508f7,
        64'h17634789_873e0367,
        64'hc783fd84_3783a6af,
        64'hf0ef853e_02c00593,
        64'h863afe44_570343dc,
        64'hfd843783_fef41223,
        64'h9be9fe44_5783fef4,
        64'h122387aa_a56ff0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_c001ae23,
        64'ha4c94785_c0e1ae23,
        64'h4705fecf_c0ef1365,
        64'h05130000_151712e5,
        64'h85930000_15972cf0,
        64'h0613a015_06f71a63,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'hc001ae23_cf91fd84,
        64'h3783fe04_1623fcf4,
        64'h2a2387ae_fca43c23,
        64'h1800f022_f4067179,
        64'h80826165_740670a6,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aaa6af_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcf984_3783baaf,
        64'hf0ef853e_02800593,
        64'h863a0ff7_7713fe44,
        64'h270343dc_f9843783,
        64'hfef42223_0047e793,
        64'hfe442783_fef42223,
        64'h87aab9cf_f0ef853e,
        64'h02800593_43dcf984,
        64'h3783ab7f_c0ef3e80,
        64'h0513a09d_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h708000ef_f9843503,
        64'h02f71163_479d873e,
        64'h57fcf984_3783a849,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_0b8000ef,
        64'hf9843503_85be5f9c,
        64'hf9843783_bc0ff0ef,
        64'h853e0300_05934609,
        64'h43dcf984_3783dfc5,
        64'h27818b89_fe442783,
        64'ha8d1fef4_26234785,
        64'hbe4ff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8f984_3783c385,
        64'h27818ff9_67a1fe44,
        64'h2703fef4_222387aa,
        64'hbd2ff0ef_853e0300,
        64'h059343dc_f9843783,
        64'haa11fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aabd8f,
        64'he0eff984_35036000,
        64'h0593863e_4681fe84,
        64'h2783df98_5007071b,
        64'h03197737_f9843783,
        64'hfef42423_1007879b,
        64'h03b907b7_a831df98,
        64'h5007071b_03197737,
        64'hf9843783_fef42423,
        64'h1007879b_03b907b7,
        64'h02f71063_4791873e,
        64'h57fcf984_3783a099,
        64'hdf982007_071b0beb,
        64'hc737f984_3783fef4,
        64'h24232007_879b03b9,
        64'h07b702f7_1063479d,
        64'h873e57fc_f9843783,
        64'ha275fef4_26234785,
        64'h14078963_2781fec4,
        64'h2783fef4_262387aa,
        64'h1d4000ef_f9843503,
        64'h50078593_031977b7,
        64'hdf985007_071b0319,
        64'h7737f984_3783ceaf,
        64'hf0ef853e_03000593,
        64'h460943dc_f9843783,
        64'hdfc52781_8b89fe44,
        64'h2783aafd_fef42623,
        64'h4785d0ef_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_f9843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aacfcf_f0ef853e,
        64'h03000593_43dcf984,
        64'h3783ac3d_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hd02fe0ef_f9843503,
        64'h60000593_863e4681,
        64'hfe842783_fef42423,
        64'h1007879b_03b907b7,
        64'h0cf71663_4789873e,
        64'h0347c783_f9843783,
        64'ha451fef4_26234785,
        64'h22078563_2781fec4,
        64'h2783fef4_262387aa,
        64'h2ac000ef_f9843503,
        64'h85be5f9c_f9843783,
        64'hdf980807_071b02fa,
        64'hf737f984_3783dc2f,
        64'hf0ef853e_03000593,
        64'h460943dc_f9843783,
        64'hdfc52781_8b89fe44,
        64'h2783acd9_fef42623,
        64'h4785de6f_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_f9843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aadd4f_f0ef853e,
        64'h03000593_43dcf984,
        64'h3783ae19_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hddafe0ef_f9843503,
        64'h60000593_863e4685,
        64'hfe842783_fef42423,
        64'h37c58100_07b7c2e1,
        64'h90234745_7010d073,
        64'h70105073_0ff0000f,
        64'h818ff0ef_f9843503,
        64'h85be863a_fa040713,
        64'h2781fe24_5783e7af,
        64'hf0ef853e_4591863a,
        64'hfe045703_43dcf984,
        64'h3783fef4_10238ff9,
        64'h17fd6785_fe045703,
        64'hfef41023_04000793,
        64'hfef41123_4785a65d,
        64'h4785c0e1_ae234705,
        64'hbf3fc0ef_53c50513,
        64'h00001517_53458593,
        64'h00001597_20400613,
        64'ha01514f7_13634785,
        64'h873e0347_c783f984,
        64'h3783c001_ae23aef9,
        64'h4785c0e1_ae234705,
        64'hc2bfc0ef_57450513,
        64'h00001517_56c58593,
        64'h00001597_20300613,
        64'ha01502f7_1f631117,
        64'h87931111_17b7873e,
        64'h53dcf984_3783c001,
        64'hae23cf91_f9843783,
        64'hfc043c23_fc043823,
        64'hfc043423_fc043023,
        64'hfa043c23_fa043823,
        64'hfa043423_fa043023,
        64'hf8a43c23_1880f0a2,
        64'hf4867159_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aaebef,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfc84,
        64'h3783f7ef_f0ef853e,
        64'h03000593_460943dc,
        64'hfc843783_dfc52781,
        64'h8b89fdc4_2783a83d,
        64'hfef42623_4785fa2f,
        64'hf0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfc843783_c3852781,
        64'h8ff967a1_fdc42703,
        64'hfcf42e23_87aaf90f,
        64'hf0ef853e_03000593,
        64'h43dcfc84_3783a8bd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_f96fe0ef,
        64'hfc843503_60000593,
        64'h863e4685_fe042783,
        64'h7010d073_70105073,
        64'h0ff0000f_fef42023,
        64'h37c10100_07b7c2e1,
        64'h90234745_9d4ff0ef,
        64'hfc843503_85befc04,
        64'h36032781_fe645783,
        64'h835ff0ef_853e4591,
        64'h863afe44_570343dc,
        64'hfc843783_fef41223,
        64'h8ff917fd_6785fe44,
        64'h5703fef4_12230400,
        64'h0793fef4_13234785,
        64'hfce7dee3_03f00793,
        64'h0007871b_fe842783,
        64'hfef42423_2785fe84,
        64'h27830007_802397ba,
        64'hfc043703_fe842783,
        64'haa154785_c0e1ae23,
        64'h4705dd5f_c0ef71e5,
        64'h05130000_15177165,
        64'h85930000_15971a80,
        64'h0613a835_fe042423,
        64'hc001ae23_a2854785,
        64'hc0e1ae23_4705e01f,
        64'hc0ef74a5_05130000,
        64'h15177425_85930000,
        64'h15971a70_0613a015,
        64'h02f71963_11178793,
        64'h111117b7_873e53dc,
        64'hfc843783_c001ae23,
        64'hcf91fc84_3783fcb4,
        64'h3023fca4_34230080,
        64'hf822fc06_71398082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'h879ff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_939ff0ef,
        64'h853e03e0_0593863a,
        64'h93411742_fe842703,
        64'h43dcfd84_3783fef4,
        64'h24238fd9_fe842783,
        64'h57f8fd84_3783fef4,
        64'h24238ff9_17e167c1,
        64'hfe842703_fef42423,
        64'h87aa93df_f0ef853e,
        64'h03e00593_43dcfd84,
        64'h378304f7_19634791,
        64'h873e57fc_fd843783,
        64'ha15ff0ef_853e0280,
        64'h0593863a_0ff77713,
        64'hfe842703_43dcfd84,
        64'h3783fef4_24230027,
        64'he793fe84_2783a039,
        64'hfef42423_0207e793,
        64'hfe842783_00f71963,
        64'h478d873e_0377c783,
        64'hfd843783_fef42423,
        64'h87aaa25f_f0ef853e,
        64'h02800593_43dcfd84,
        64'h378393ef_d0ef3e80,
        64'h05139f7f_f0ef853e,
        64'h03000593_460943dc,
        64'hfd843783_dfc52781,
        64'h8b89fe84_2783a8f5,
        64'hfef42623_4785a1bf,
        64'hf0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c3852781,
        64'h8ff967a1_fe842703,
        64'hfef42423_87aaa09f,
        64'hf0ef853e_03000593,
        64'h43dcfd84_3783aa35,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_a0ffe0ef,
        64'hfd843503_60000593,
        64'h863e4681_fe442783,
        64'hfef42223_1007879b,
        64'h03b707b7_a039fef4,
        64'h22235007_879b03b7,
        64'h07b700f7_19634791,
        64'h873e57fc_fd843783,
        64'ha02dfef4_22232007,
        64'h879b03b7_07b7a825,
        64'hfef42223_6007879b,
        64'h03b707b7_00f71963,
        64'h4791873e_57fcfd84,
        64'h378302f7_1763478d,
        64'h873e0377_c783fd84,
        64'h378302e7_8ba34709,
        64'hfd843783_a03102e7,
        64'h8ba3470d_fd843783,
        64'h00f71863_47a1873e,
        64'h4bdcfd84_378300f7,
        64'h1f634795_873e0347,
        64'hc783fd84_378302f7,
        64'h17634789_873e0367,
        64'hc783fd84_3783a431,
        64'hfef42623_47851207,
        64'h8c632781_fec42783,
        64'hfef42623_87aaae1f,
        64'he0effd84_35036007,
        64'h859367a1_863e4681,
        64'hfe442783_fef42223,
        64'h0377c783_fd843783,
        64'h02e78ba3_4709fd84,
        64'h3783ac81_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hb23fe0ef_fd843503,
        64'h70078593_678d863e,
        64'h46814bbc_fd843783,
        64'h06f71b63_4785873e,
        64'h0347c783_fd843783,
        64'ha479fe04_262300e7,
        64'he563478d_873e4bdc,
        64'hfd843783_a45d4785,
        64'hc0e1ae23_4705900f,
        64'hd0efa4a5_05130000,
        64'h2517a425_85930000,
        64'h259711b0_0613a015,
        64'h02f71e63_4789873e,
        64'h0367c783_fd843783,
        64'hc001ae23_acf94785,
        64'hc0e1ae23_4705938f,
        64'hd0efa825_05130000,
        64'h2517a7a5_85930000,
        64'h259711a0_0613a015,
        64'h02f71f63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_c001ae23,
        64'hcf91fd84_3783fca4,
        64'h3c231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_badff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fd843783,
        64'hc6dff0ef_853e0300,
        64'h05934609_43dcfd84,
        64'h3783dfc5_27818b89,
        64'hfe042783_a83dfef4,
        64'h26234785_c91ff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c385_27818ff9,
        64'h67a1fe04_2703fef4,
        64'h202387aa_c7fff0ef,
        64'h853e0300_059343dc,
        64'hfd843783_a8bdfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aac85f_e0effd84,
        64'h35033007_859367ad,
        64'h460186be_2781fe64,
        64'h57837010_d0737010,
        64'h50730ff0_000fc2e1,
        64'h90234745_ebcff0ef,
        64'hfd843503_85befd04,
        64'h36032781_fe645783,
        64'hd1dff0ef_853e4591,
        64'h863afe44_570343dc,
        64'hfd843783_fef41223,
        64'h8ff917fd_6785fe44,
        64'h5703fef4_122347a1,
        64'hfef41323_4785a201,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_d07fe0ef,
        64'hfd843503_70078593,
        64'h678d863e_46814bbc,
        64'hfd843783_fce7dfe3,
        64'h479d0007_871bfe84,
        64'h2783fef4_24232785,
        64'hfe842783_00078023,
        64'h97bafd04_3703fe84,
        64'h2783aaa1_4785c0e1,
        64'hae234705_ae6fd0ef,
        64'hc3050513_00002517,
        64'hc2858593_00002597,
        64'h0ba00613_a835fe04,
        64'h2423c001_ae23a251,
        64'h4785c0e1_ae234705,
        64'hb12fd0ef_c5c50513,
        64'h00002517_c5458593,
        64'h00002597_0b900613,
        64'ha01502f7_19631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783c001,
        64'hae23cf91_fd843783,
        64'hfcb43823_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623e2ff_f0ef8536,
        64'h4591863e_93c117c2,
        64'h8ff917fd_6785fd64,
        64'h570343d4_fd843783,
        64'hfef42623_278187aa,
        64'hda9ff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_a081fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aae25f_e0effd84,
        64'h35036585_863e4681,
        64'h2781fd64_5783a0ad,
        64'hfef42623_4785a89d,
        64'h4785c0e1_ae234705,
        64'hbe2fd0ef_d2c50513,
        64'h00002517_d2458593,
        64'h00002597_07f00613,
        64'ha015c79d_27813037,
        64'hf793fe84_2783fef4,
        64'h242387aa_e25ff0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783c001_ae23a0d9,
        64'h4785c0e1_ae234705,
        64'hc32fd0ef_d7c50513,
        64'h00002517_d7458593,
        64'h00002597_07e00613,
        64'ha01504f7_1b631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783c001,
        64'hae23cf91_fd843783,
        64'hfcf41b23_87aefca4,
        64'h3c231800_f022f406,
        64'h71798082_61056442,
        64'h60e20001_eb7ff0ef,
        64'h853e85ba_fea44703,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_052387ba,
        64'hfef405a3_87b6fef4,
        64'h26238732_86ae87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h853e87aa_ea9ff0ef,
        64'h853e9381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef405a3,
        64'h87bafef4_2623872e,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e20001_f63ff0ef,
        64'h853e85ba_fe845703,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_142387ba,
        64'hfef405a3_87b6fef4,
        64'h26238732_86ae87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h853e87aa_f47ff0ef,
        64'h853e9381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef405a3,
        64'h87bafef4_2623872e,
        64'h87aa1000_e822ec06,
        64'h11018082_61457422,
        64'h000100e7_9023fd64,
        64'h5703fe84_3783fef4,
        64'h3423fd84_3783fcf4,
        64'h1b2387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61457422_000100e7,
        64'h8023fd74_4703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_0ba387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61056462,
        64'h853e2781_439cfe84,
        64'h3783fea4_34231000,
        64'hec221101_80826105,
        64'h6462853e_93c117c2,
        64'h0007d783_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61056462,
        64'h853e0ff7_f7930007,
        64'hc783fe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826161_640660a6,
        64'h853efec4_2783fe04,
        64'h2623d3f8_fb843783,
        64'h0007871b_0097d79b,
        64'hfd842783_fcf42c23,
        64'h02f707bb_fe042783,
        64'hfd842703_fcf42c23,
        64'h02f707bb_fdc42703,
        64'h27812785_fd842783,
        64'hfcf42c23_8fd9fd84,
        64'h27830007_871b8ff9,
        64'hc0078793_6785873e,
        64'h278100a7_979bfd04,
        64'h2783fcf4_2c230167,
        64'hd79bfcc4_2783fcf4,
        64'h2e232781_00f717bb,
        64'h47052781_27892781,
        64'h8b9d2781_0077d79b,
        64'hfcc42783_fef42023,
        64'h278100f7_17bb4705,
        64'h27818bbd_27810087,
        64'hd79bfd04_278302e7,
        64'h8aa3fb84_37830ff7,
        64'hf7138bbd_0ff7f793,
        64'h27810127_d79bfd44,
        64'h2783fcf4_2a232781,
        64'h87aaa11f_d0ef853e,
        64'h93811782_278127f1,
        64'h43dcfb84_3783fcf4,
        64'h28232781_87aaa2df,
        64'hd0ef853e_93811782,
        64'h278127e1_43dcfb84,
        64'h3783fcf4_26232781,
        64'h87aaa49f_d0ef853e,
        64'h93811782_278127d1,
        64'h43dcfb84_3783fcf4,
        64'h24232781_87aaa65f,
        64'hd0ef853e_93811782,
        64'h278127c1_43dcfb84,
        64'h3783a23d_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h9e2ff0ef_fb843503,
        64'h90078593_6785863e,
        64'h46814bbc_fb843783,
        64'haab1fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaa10f,
        64'hf0effb84_35033000,
        64'h0593863e_46814bbc,
        64'hfb843783_cbb81234,
        64'h0737fb84_3783c7f8,
        64'hfb843783_0007871b,
        64'h87aab85f_d0ef853e,
        64'h45f143dc_fb843783,
        64'hc7b8fb84_37830007,
        64'h871b87aa_b9ffd0ef,
        64'h853e45e1_43dcfb84,
        64'h3783c3f8_fb843783,
        64'h0007871b_87aabb9f,
        64'hd0ef853e_45d143dc,
        64'hfb843783_c3b8fb84,
        64'h37830007_871b87aa,
        64'hbd3fd0ef_853e45c1,
        64'h43dcfb84_3783aaed,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_aaeff0ef,
        64'hfb843503_20000593,
        64'h46014681_db984705,
        64'hfb843783_c7892781,
        64'h8ff94000_07b7fe84,
        64'h2703fa07_dde3fe84,
        64'h2783fef4_242387aa,
        64'hb8ffd0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_aca1fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aab0cf_f0effb84,
        64'h35031000_059340ff,
        64'h86374681_a091fe04,
        64'h2423a459_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hb3aff0ef_fb843503,
        64'h45814601_4681a46d,
        64'hfef42623_4785e789,
        64'h27818ff9_67c1fe44,
        64'h2703fef4_222387aa,
        64'hc0ffd0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfb84_3783cb8d,
        64'h47dcfb84_378302f7,
        64'h0e634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_fb843783,
        64'ha6014785_c0e1ae23,
        64'h470593df_d0ef2665,
        64'h05130000_25172665,
        64'h85930000_25976890,
        64'h0613a015_04f71163,
        64'h4789873e_0367c783,
        64'hfb843783_c001ae23,
        64'hae254785_c0e1ae23,
        64'h4705975f_d0ef29e5,
        64'h05130000_251729e5,
        64'h85930000_25976880,
        64'h0613a015_02f71f63,
        64'h11178793_111117b7,
        64'h873e53dc_fb843783,
        64'hc001ae23_cf91fb84,
        64'h3783faa4_3c230880,
        64'he0a2e486_715d8082,
        64'h61217442_70e20001,
        64'h7010d073_70105073,
        64'h0ff0000f_d55fd0ef,
        64'h853a85be_27810807,
        64'h8793fd84_37839301,
        64'h02079713_27810587,
        64'h879b43dc_fd843783,
        64'h00e79123_97b6078e,
        64'h07c19381_02061793,
        64'hfd843683_93410307,
        64'h971302f7_07bb0006,
        64'h861b36fd_fec42683,
        64'h93c117c2_fe442783,
        64'h93410307_9713fd44,
        64'h278300e7_90230230,
        64'h071397ba_078e07c1,
        64'h93811782_fd843703,
        64'h278137fd_fec42783,
        64'hc3d897b6_078e07c1,
        64'h93810206_1793fd84,
        64'h36830007_871b9fb9,
        64'h0006861b_36fdfec4,
        64'h26832781_0107979b,
        64'hfe842783_0007871b,
        64'hfc843783_f8e7ebe3,
        64'h2781fe84_27830007,
        64'h871b37fd_fec42783,
        64'hfef42423_2785fe84,
        64'h27830007_912397ba,
        64'h078e07c1_fe846783,
        64'hfd843703_00e79023,
        64'h02100713_97ba078e,
        64'h07c1fe84_6783fd84,
        64'h3703c3d8_97b6078e,
        64'h07c1fe84_6783fd84,
        64'h36830007_871b9fb9,
        64'h27810107_979bfe84,
        64'h27830007_871bfc84,
        64'h3783a8b1_fe042423,
        64'hfef42623_2785fec4,
        64'h2783c791_27818ff9,
        64'h17fd67c1_873e2781,
        64'h02f707bb_fe442783,
        64'hfd442703_fef42623,
        64'h0107d79b_278102f7,
        64'h07bbfe44_2783fd44,
        64'h2703a835_fef42623,
        64'h478500f7_766367c1,
        64'h873e2781_02f707bb,
        64'hfe442783_fd442703,
        64'hfef42223_8ff917fd,
        64'h6785fe44_2703fef4,
        64'h222387aa_f0ffd0ef,
        64'h853e4591_43dcfd84,
        64'h3783fe04_2223fe04,
        64'h2423fe04_2623fcf4,
        64'h2a23fcc4_342387ae,
        64'hfca43c23_0080f822,
        64'hfc067139_80826145,
        64'h740270a2_853efec4,
        64'h27830001_a011fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aae1cf_f0effd84,
        64'h35037000_0593863e,
        64'h46814bbc_fd843783,
        64'hfe042623_fca43c23,
        64'h1800f022_f4067179,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623fd7f_d0ef853e,
        64'h03000593_460943dc,
        64'hfd843783_dfc52781,
        64'h8b89fe44_2783a00d,
        64'hfef42623_4785ffbf,
        64'hd0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c3852781,
        64'h8ff967a1_fe442703,
        64'hfef42223_87aafe9f,
        64'hd0ef853e_03000593,
        64'h43dcfd84_3783a08d,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_ec6ff0ef,
        64'hfd843503_90078593,
        64'h6789863e_86bafd44,
        64'h2783fd04_2703c2e1,
        64'h90230270_0713a869,
        64'hfef42623_4785c3a9,
        64'h2781fec4_2783fef4,
        64'h262387aa_efeff0ef,
        64'hfd843503_80078593,
        64'h6789863e_86bafd44,
        64'h2783fd04_2703c2e1,
        64'h9023470d_02f71d63,
        64'h47850007_871bfd04,
        64'h27837010_d0737010,
        64'h50730ff0_000f1460,
        64'h00effd84_350385be,
        64'hfc843603_fd042783,
        64'ha8f5fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa0810,
        64'h00effd84_35032000,
        64'h059302f7_03632000,
        64'h0793873e_278187aa,
        64'h826fe0ef_853e9381,
        64'h17822781_279143dc,
        64'hfd843783_a281fef4,
        64'h26234785_e7892781,
        64'h8ff967c1_fe842703,
        64'hfef42423_87aa854f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_cb8d47dc,
        64'hfd843783_02f70e63,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cfd84_378300f7,
        64'h1f634789_873e0367,
        64'hc783fd84_3783fcf4,
        64'h282387ba_fcf42a23,
        64'hfcd43423_873287ae,
        64'hfca43c23_0080f822,
        64'hfc067139_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aa8d4f,
        64'he0ef853e_93811782,
        64'h278127c1_43dcfd84,
        64'h37839bef_e0ef853e,
        64'h03000593_460943dc,
        64'hfd843783_dfc52781,
        64'h8b89fe44_2783a83d,
        64'hfef42623_47859e2f,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c3852781,
        64'h8ff967a1_fe442703,
        64'hfef42223_87aa9d0f,
        64'he0ef853e_03000593,
        64'h43dcfd84_3783a8bd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_8afff0ef,
        64'hfd843503_20078593,
        64'h6785863e_86bafd44,
        64'h2783fd04_2703c2e1,
        64'h90230370_0713a85d,
        64'hfef42623_4785c3a9,
        64'h2781fec4_2783fef4,
        64'h262387aa_8e7ff0ef,
        64'hfd843503_10078593,
        64'h6785863e_86bafd44,
        64'h2783fd04_2703c2e1,
        64'h9023474d_02f71d63,
        64'h47850007_871bfd04,
        64'h27837010_d0737010,
        64'h50730ff0_000f32e0,
        64'h00effd84_350385be,
        64'hfc843603_fd042783,
        64'haa21fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa2690,
        64'h00effd84_35032000,
        64'h059302f7_03632000,
        64'h0793873e_278187aa,
        64'ha0efe0ef_853e9381,
        64'h17822781_279143dc,
        64'hfd843783_aab1fef4,
        64'h26234785_e7892781,
        64'h8ff967c1_fe842703,
        64'hfef42423_87aaa3cf,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_cb8d47dc,
        64'hfd843783_02f70e63,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cfd84_378300f7,
        64'h1f634789_873e0367,
        64'hc783fd84_3783fcf4,
        64'h282387ba_fcf42a23,
        64'hfcd43423_873287ae,
        64'hfca43c23_0080f822,
        64'hfc067139_80826145,
        64'h7422853e_fec42783,
        64'h0001a011_0001a021,
        64'h0001a031_fef42623,
        64'h8fd9fd44_2783fec4,
        64'h2703a831_fef42623,
        64'h01a7e793_fec42783,
        64'ha02dfef4_262303a7,
        64'he793fec4_2783a825,
        64'hfef42623_01a7e793,
        64'hfec42783_a099fef4,
        64'h26230027_e793fec4,
        64'h2783a891_fef42623,
        64'h03a7e793_fec42783,
        64'ha08dfef4_262303a7,
        64'he793fec4_2783a885,
        64'hfef42623_01a7e793,
        64'hfec42783_a8bdfef4,
        64'h26230097_e793fec4,
        64'h2783a071_fef42623,
        64'h03a7e793_fec42783,
        64'ha869fef4_262301a7,
        64'he793fec4_278300f7,
        64'h19634785_873e0347,
        64'hc783fd84_3783a865,
        64'hfef42623_01a7e793,
        64'hfec42783_a0d9fef4,
        64'h262301a7_e793fec4,
        64'h2783a8d1_fef42623,
        64'h01b7e793_fec42783,
        64'ha0cdfef4_262303a7,
        64'he793fec4_278300f7,
        64'h19634785_873e0347,
        64'hc783fd84_3783a201,
        64'hfef42623_01b7e793,
        64'hfec42783_a239fef4,
        64'h262301b7_e793fec4,
        64'h2783aa31_fef42623,
        64'h0097e793_fec42783,
        64'ha22dfef4_26230027,
        64'he793fec4_2783aa39,
        64'h0ef70563_90078793,
        64'h67ad0007_871b10e6,
        64'h8a633007_0713672d,
        64'h0007869b_10e68a63,
        64'ha0070713_672d0007,
        64'h869ba2a9_16f70363,
        64'ha0078793_67910007,
        64'h871b0ee6_8d63d007,
        64'h07136725_0007869b,
        64'h0ae68963_60070713,
        64'h67210007_869b02d7,
        64'h68637007_07136725,
        64'h0007869b_14e68063,
        64'h70070713_67250007,
        64'h869baa49_14f70863,
        64'h80078793_67890007,
        64'h871b18e6_8b634007,
        64'h0713670d_0007869b,
        64'h16e68663_90070713,
        64'h67090007_869baa7d,
        64'h16f70763_20078793,
        64'h67850007_871b16e6,
        64'h8e635007_07136705,
        64'h0007869b_18e68563,
        64'h30070713_67050007,
        64'h869b02d7_68637007,
        64'h07136705_0007869b,
        64'h1ae68a63_70070713,
        64'h67050007_869b06d7,
        64'h6c637007_0713670d,
        64'h0007869b_20e68463,
        64'h70070713_670d0007,
        64'h869ba40d_1cf70263,
        64'hb0078793_67850007,
        64'h871b1ce6_89636705,
        64'h0007869b_1ce68e63,
        64'hc0070713_67050007,
        64'h869ba4a9_1af70263,
        64'h70000793_0007871b,
        64'h1ee68563_90070713,
        64'h67050007_869b1c07,
        64'h06632701_8007871b,
        64'h02d76563_a0070713,
        64'h67050007_869b20e6,
        64'h8f63a007_07136705,
        64'h0007869b_a47118f7,
        64'h08633000_07930007,
        64'h871b1ae6_85635000,
        64'h07130007_869b2ae6,
        64'h8e634000_07130007,
        64'h869bac4d_18f70d63,
        64'h10000793_0007871b,
        64'h2c070963_0007871b,
        64'h00d76d63_20000713,
        64'h0007869b_1ce68463,
        64'h20000713_0007869b,
        64'h04d76c63_60000713,
        64'h0007869b_20e68563,
        64'h60000713_0007869b,
        64'h0cd76d63_10070713,
        64'h67050007_869b2ae6,
        64'h8a631007_07136705,
        64'h0007869b_fd442783,
        64'hfef42623_fd442783,
        64'hfcf42a23_87aefca4,
        64'h3c231800_f4227179,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623edef_e0ef853e,
        64'h03000593_460543dc,
        64'hfd843783_d3a92781,
        64'h8b85fe04_2783a00d,
        64'hefcfe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783fef4,
        64'h26234789_e7812781,
        64'h9bf9fec4_2783fef4,
        64'h262387aa_eeefe0ef,
        64'h853e0320_059343dc,
        64'hfd843783_c3a12781,
        64'h8ff967a1_fe042703,
        64'ha899f46f_e0ef853e,
        64'h03000593_02000613,
        64'h43dcfd84_3783cf81,
        64'h27810207_f7932781,
        64'h87aaf2cf_e0ef853e,
        64'h03000593_43dcfd84,
        64'h378302f7_1b633007,
        64'h87936785_0007871b,
        64'hfd442783_00f70b63,
        64'h50078793_67850007,
        64'h871bfd44_2783fef4,
        64'h202387aa_f66fe0ef,
        64'h853e0300_059343dc,
        64'hfd843783_f4cfe0ef,
        64'h853a85be_27818fd5,
        64'h2781c201_d7830007,
        64'h869b0107_979bfe44,
        64'h27839301_02079713,
        64'h278127b1_43dcfd84,
        64'h3783a219_fef42623,
        64'h4785c789_27810207,
        64'hf793fe44_2783cb99,
        64'h27818b89_fe842783,
        64'hfef42423_87aaf2cf,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_02f70f63,
        64'h30078793_67850007,
        64'h871bfd44_278304f7,
        64'h08635007_87936785,
        64'h0007871b_fd442783,
        64'hfef42223_8ff917fd,
        64'h6791fe44_2703fef4,
        64'h222387aa_188000ef,
        64'hfd843503_85befd44,
        64'h278385ff_e0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'h875fe0ef_853a0300,
        64'h0593fff7_861367c1,
        64'h43d8fd84_3783827f,
        64'he0ef853e_85bafd04,
        64'h27039381_17822781,
        64'h27a143dc_fd843783,
        64'h925fe0ef_853e02e0,
        64'h05934639_43dcfd84,
        64'h37838b7f_e0ef853e,
        64'h4599863a_93411742,
        64'hfcc42703_43dcfd84,
        64'h3783aadd_fef42623,
        64'h4785a409_4785c0e1,
        64'hae234705_cf6fe0ef,
        64'he2050513_00003517,
        64'he2058593_00003597,
        64'h44c00613_a015c79d,
        64'h27818b85_fe842783,
        64'hfef42423_87aa835f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_c001ae23,
        64'hac814785_c0e1ae23,
        64'h4705d44f_e0efe6e5,
        64'h05130000_3517e6e5,
        64'h85930000_359744b0,
        64'h0613a015_04f71a63,
        64'h11178793_111117b7,
        64'h873e53dc_fd843783,
        64'hc001ae23_cf91fd84,
        64'h3783fcf4_262387ba,
        64'hfcf42823_87b2fcf4,
        64'h2a238736_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_61457402,
        64'h70a2853e_fec42783,
        64'h0001fcf7_19e301f0,
        64'h07b7873e_27818ff9,
        64'h01f007b7_fe842703,
        64'hfef42423_87aa8ddf,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_a839fef4,
        64'h242387aa_8fbfe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h378380ff_e0ef3e80,
        64'h05139eff_e0ef853a,
        64'h02c00593_863e93c1,
        64'h17c20047_e79393c1,
        64'h17c2fe44_278343d8,
        64'hfd843783_fef42223,
        64'h87aa9ddf_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783d3ed_27818b89,
        64'hfe442783_fef42223,
        64'h87aa9fdf_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783a821_fef42223,
        64'h87aaa15f_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783a5ff_e0ef853a,
        64'h02c00593_863e93c1,
        64'h17c20017_e79393c1,
        64'h17c2fe44_278343d8,
        64'hfd843783_fef42223,
        64'h87aaa4df_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783a211_fef42623,
        64'h4785e789_27818ba1,
        64'h2781fe24_5783fef4,
        64'h112387aa_a77fe0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_8e9fe0ef,
        64'h38878513_6785acbf,
        64'he0ef853e_03e00593,
        64'h863afe24_570343dc,
        64'hfd843783_fef41123,
        64'h0087e793_fe245783,
        64'hfef41123_87aaab9f,
        64'he0ef853e_03e00593,
        64'h43dcfd84_3783b03f,
        64'he0ef853e_02c00593,
        64'h863afe24_570343dc,
        64'hfd843783_fef41123,
        64'h9be9fe24_5783fef4,
        64'h112387aa_aeffe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_ffe12781,
        64'h8ff901f0_07b7fe84,
        64'h2703fef4_242387aa,
        64'ha77fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783a839,
        64'hfef42423_87aaa95f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_fef42623,
        64'h4785c781_2781fec4,
        64'h2783fef4_262387aa,
        64'h212000ef_fd843503,
        64'hb0078593_67854601,
        64'h4681fca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'hf3e52781_8b892781,
        64'hfeb44783_fef405a3,
        64'h87aac1df_e0ef853e,
        64'h02f00593_43dcfd84,
        64'h3783a821_fef405a3,
        64'h87aac35f_e0ef853e,
        64'h02f00593_43dcfd84,
        64'h3783c7ff_e0ef853e,
        64'h02f00593_460943dc,
        64'hfd843783_c11fe0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c27f_e0ef853a,
        64'h03000593_fff78613,
        64'h67c143d8_fd843783,
        64'h02e78a23_4709fd84,
        64'h3783a031_02e78a23,
        64'h4705fd84_3783c799,
        64'h2781fec4_2783fef4,
        64'h262387aa_2de000ef,
        64'hfd843503_10000593,
        64'h40ff8637_4681a855,
        64'hfef42623_4785a0c1,
        64'h4785c0e1_ae234705,
        64'h89bfe0ef_1c450513,
        64'h00003517_1c458593,
        64'h00003597_3ac00613,
        64'ha015c79d_2781fec4,
        64'h2783fef4_262387aa,
        64'h32a000ef_fd843503,
        64'h45814601_4681ae3f,
        64'he0ef7107_85136789,
        64'hc001ae23_a2394785,
        64'hc0e1ae23_47058e9f,
        64'he0ef2125_05130000,
        64'h35172125_85930000,
        64'h35973ab0_0613a015,
        64'h04f71a63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_c001ae23,
        64'hcf91fd84_3783fca4,
        64'h3c231800_f022f406,
        64'h71798082_614d64ea,
        64'h740a70aa_853efdc4,
        64'h27830001_a0110001,
        64'ha0210001_a031fcf4,
        64'h2e234785_cb892781,
        64'hfdc42783_fcf42e23,
        64'h87aa4e40_10eff584,
        64'h35032000_059302f7,
        64'h17634785_873e0347,
        64'hc783f584_378300f7,
        64'h1a634791_873e57fc,
        64'hf5843783_0001a0b9,
        64'hfcf42e23_4785c791,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_71e020ef,
        64'hf5843503_85befd44,
        64'h2783fcf4_2a231007,
        64'h879b03a2_07b7eb95,
        64'h0a27c783_6b478793,
        64'h1ffed797_a071fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa0650_10eff584,
        64'h350302f7_11634791,
        64'h873e57fc_f5843783,
        64'ha865fcf4_2e234785,
        64'h00f70663_4785873e,
        64'h0b97c783_6fc78793,
        64'h1ffed797_04f71663,
        64'h4791873e_57fcf584,
        64'h378300f7_09634795,
        64'h873e57fc_f5843783,
        64'ha8c5fcf4_2e234785,
        64'h00f70663_4789873e,
        64'h0b97c783_73478793,
        64'h1ffed797_02f71063,
        64'h479d873e_57fcf584,
        64'h3783aa29_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h634020ef_f5843503,
        64'h76858593_1ffed597,
        64'ha281fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa6070,
        64'h10eff584_35030cf7,
        64'h0b634799_873e57fc,
        64'hf5843783_d7f84719,
        64'hf5843783_a029d7f8,
        64'h4715f584_378300e7,
        64'hf7634785_873e0377,
        64'hc783f584_3783cf91,
        64'h27818b89_27810c47,
        64'hc7837ca7_87931ffe,
        64'hd797a825_d7f84711,
        64'hf5843783_00e7f763,
        64'h4785873e_0377c783,
        64'hf5843783_cf912781,
        64'h8bb12781_0c47c783,
        64'h7f878793_1ffed797,
        64'ha09dd7f8_471df584,
        64'h378300e7_f7634785,
        64'h873e0377_c783f584,
        64'h3783cf91_27810307,
        64'hf7932781_0c47c783,
        64'h82878793_1ffee797,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810d47,
        64'hc7838427_87931ffe,
        64'he79753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810087,
        64'h979b2781_0d57c783,
        64'h86878793_1ffee797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h8fd92781_0107979b,
        64'h27810d67_c78388e7,
        64'h87931ffe_e79753f8,
        64'hf5843783_d3f8f584,
        64'h37830007_871b0187,
        64'h979b2781_0d77c783,
        64'h8b078793_1ffee797,
        64'ha461fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa7a20,
        64'h20eff584_35038d65,
        64'h85931ffe_e597a47d,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_287010ef,
        64'hf5843503_28f71263,
        64'h4795873e_0347c783,
        64'hf5843783_acf1fcf4,
        64'h2e234785_28f70d63,
        64'h4785873e_0b97c783,
        64'h92078793_1ffee797,
        64'hace5fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa0130,
        64'h20eff584_35039465,
        64'h85931ffe_e597ae39,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_7e5010ef,
        64'hf5843503_d7f84715,
        64'hf5843783_2ee7fd63,
        64'h4785873e_0377c783,
        64'hf5843783_30078563,
        64'h27818b89_27810c47,
        64'hc7839927_87931ffe,
        64'he797d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0d47c783_9ac78793,
        64'h1ffee797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0087979b_27810d57,
        64'hc7839d27_87931ffe,
        64'he79753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810107,
        64'h979b2781_0d67c783,
        64'h9f878793_1ffee797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h0187979b_27810d77,
        64'hc783a1a7_87931ffe,
        64'he797aecd_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h10d020ef_f5843503,
        64'ha4058593_1ffee597,
        64'ha921fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa3f10,
        64'h10eff584_350314f7,
        64'h1f634785_873e0367,
        64'hc783f584_378316e7,
        64'hf763478d_873e0357,
        64'hc783f584_378316f7,
        64'h1f634789_873e0347,
        64'hc783f584_3783a19d,
        64'hfcf42e23_47854207,
        64'h83632781_fdc42783,
        64'hfcf42e23_87aa12e0,
        64'h20eff584_3503d7f8,
        64'h4715f584_378344e7,
        64'hf3634785_873e0377,
        64'hc783f584_37834407,
        64'h8b632781_8b892781,
        64'hf9d44783_46078263,
        64'h0004c783_02e78e23,
        64'h4705f584_378380af,
        64'hf0ef3e80_05139eaf,
        64'hf0ef853a_02c00593,
        64'h863e93c1_17c20047,
        64'he793fda4_578343d8,
        64'hf5843783_fcf41d23,
        64'h87aa9d4f_f0ef853e,
        64'h02c00593_43dcf584,
        64'h3783d3e5_27818b89,
        64'h2781fda4_5783fcf4,
        64'h1d2387aa_9f6ff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_a821fcf4,
        64'h1d2387aa_a0eff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_a58ff0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0017e793,
        64'hfda45783_43d8f584,
        64'h3783fcf4_1d2387aa,
        64'ha42ff0ef_853e02c0,
        64'h059343dc_f5843783,
        64'ha3a5fcf4_2e234785,
        64'he7892781_8ba12781,
        64'hfd245783_fcf41923,
        64'h87aaa6cf_f0ef853e,
        64'h03e00593_43dcf584,
        64'h37838def_f0ef3887,
        64'h85136785_ac0ff0ef,
        64'h853e03e0_0593863a,
        64'hfd245703_43dcf584,
        64'h3783fcf4_19230087,
        64'he793fd24_5783fcf4,
        64'h192387aa_aaeff0ef,
        64'h853e03e0_059343dc,
        64'hf5843783_af8ff0ef,
        64'h853e02c0_0593863a,
        64'hfd245703_43dcf584,
        64'h3783fcf4_19239be9,
        64'hfd245783_fcf41923,
        64'h87aaae4f_f0ef853e,
        64'h02c00593_43dcf584,
        64'h37831407_9d6303c7,
        64'hc783f584_378316f7,
        64'h136347a1_873e4bdc,
        64'hf5843783_16e7fa63,
        64'h478d873e_f9d44783,
        64'h1807d063_4187d79b,
        64'h0187979b_0024c783,
        64'h62079e63_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h146020ef_f5843503,
        64'h85bef904_0793adb9,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_637010ef,
        64'hf5843503_c3852781,
        64'h8b912781_0014c783,
        64'ha561fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa4830,
        64'h10eff584_350385a6,
        64'ha565fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa2e50,
        64'h20eff584_350326f7,
        64'h12634785_873e0347,
        64'hc783f584_3783add9,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_450010ef,
        64'hf5843503_add5fcf4,
        64'h2e234785_adf5fcf4,
        64'h2e234785_cb892781,
        64'hfdc42783_fcf42e23,
        64'h87aa0170_20eff584,
        64'h350385be_5f9cf584,
        64'h3783df98_a807071b,
        64'h018cc737_f5843783,
        64'haf05fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa6cc0,
        64'h10eff584_350304f7,
        64'h1b634795_873e0347,
        64'hc783f584_378300f7,
        64'h0a634789_873e0347,
        64'hc783f584_3783a7bd,
        64'hfcf42e23_4785c3d1,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_089020ef,
        64'hf5843503_85be5f9c,
        64'hf5843783_df988407,
        64'h071b017d_8737f584,
        64'h3783a801_df98ac07,
        64'h071b0121_f737f584,
        64'h378300f7_1a634789,
        64'h873e0367_c783f584,
        64'h37837c40_006ffcf4,
        64'h2e234785_c7912781,
        64'hfdc42783_fcf42e23,
        64'h87aa935f_f0eff584,
        64'h350306f7_1c634785,
        64'h873e0347_c783f584,
        64'h37837f40_006ffcf4,
        64'h2e234785_00f70763,
        64'h4795873e_0347c783,
        64'hf5843783_00f70f63,
        64'h4789873e_0347c783,
        64'hf5843783_02f70763,
        64'h4785873e_0347c783,
        64'hf5843783_02f702e3,
        64'h47850007_871bfdc4,
        64'h2783fcf4_2e2387aa,
        64'h053000ef_f5843503,
        64'ha83902e7_8a234715,
        64'hf5843783_00f71863,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cf584_37830750,
        64'h006f4785_c0e1ae23,
        64'h47059b4f_f0efade5,
        64'h05130000_4517ade5,
        64'h85930000_45972400,
        64'h0613a01d_04f71863,
        64'h4789873e_0367c783,
        64'hf5843783_df98a807,
        64'h071b0006_2737f584,
        64'h37830207_8e23f584,
        64'h378302e7_8a234705,
        64'hf5843783_02e78ba3,
        64'h4705f584_3783c001,
        64'hae230d90_006f4785,
        64'hc0e1ae23_4705a18f,
        64'hf0efb425_05130000,
        64'h4517b425_85930000,
        64'h459723f0_0613a01d,
        64'h06f71563_11178793,
        64'h111117b7_873e53dc,
        64'hf5843783_c001ae23,
        64'hcf91f584_3783fc04,
        64'h3423fc04_3023fa04,
        64'h3c23fa04_3823fa04,
        64'h3423fa04_3023f804,
        64'h3c23f804_38230004,
        64'hb0230057_94938395,
        64'h07fdf807_8793fe04,
        64'h0793f4a4_3c231900,
        64'hed26f122_f5067171,
        64'h80826161_640660a6,
        64'h853efec4_2783fe04,
        64'h2623d3f8_fb843783,
        64'h0007871b_00a7979b,
        64'h27812785_27818ff9,
        64'h17fd0040_07b7873e,
        64'h27810087_d79bfc44,
        64'h278302f7_16634785,
        64'h873e2781_8b8d2781,
        64'h0167d79b_fcc42783,
        64'ha081d3f8_fb843783,
        64'h0007871b_0097d79b,
        64'hfd042783_fcf42823,
        64'h02f707bb_fd842783,
        64'hfd042703_fcf42823,
        64'h02f707bb_fd442703,
        64'h27812785_fd042783,
        64'hfcf42823_8fd9fd04,
        64'h27830007_871b8ff9,
        64'hc0078793_6785873e,
        64'h278100a7_979bfc84,
        64'h2783fcf4_28230167,
        64'hd79bfc44_2783fcf4,
        64'h2a232781_00f717bb,
        64'h47052781_27892781,
        64'h8b9d2781_0077d79b,
        64'hfc442783_fcf42c23,
        64'h278100f7_17bb4705,
        64'h27818bbd_27810087,
        64'hd79bfc84_2783e3c5,
        64'h27818b8d_27810167,
        64'hd79bfcc4_2783fcf4,
        64'h26232781_87aaeacf,
        64'hf0ef853e_93811782,
        64'h278127f1_43dcfb84,
        64'h3783fcf4_24232781,
        64'h87aaec8f_f0ef853e,
        64'h93811782_278127e1,
        64'h43dcfb84_3783fcf4,
        64'h22232781_87aaee4f,
        64'hf0ef853e_93811782,
        64'h278127d1_43dcfb84,
        64'h3783fcf4_20232781,
        64'h87aaf00f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783a28d,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_67f000ef,
        64'hfb843503_90078593,
        64'h6785863e_46814bbc,
        64'hfb843783_d7d54bbc,
        64'hfb843783_cbb8fb84,
        64'h37830007_871b8ff9,
        64'h77c1873e_278187aa,
        64'hf5eff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_a2c1fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa6dd0_00effb84,
        64'h35033000_05934601,
        64'h4681c7f8_fb843783,
        64'h0007871b_87aa841f,
        64'hf0ef853e_45f143dc,
        64'hfb843783_c7b8fb84,
        64'h37830007_871b87aa,
        64'h85bff0ef_853e45e1,
        64'h43dcfb84_3783c3f8,
        64'hfb843783_0007871b,
        64'h87aa875f_f0ef853e,
        64'h45d143dc_fb843783,
        64'hc3b8fb84_37830007,
        64'h871b87aa_88fff0ef,
        64'h853e45c1_43dcfb84,
        64'h3783a4b9_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h76b000ef_fb843503,
        64'h20000593_46014681,
        64'hac95fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa5650,
        64'h00effb84_350302e7,
        64'h8e234705_fb843783,
        64'hc78d2781_8ff90100,
        64'h07b7fe84_2703db98,
        64'h4705fb84_3783c789,
        64'h27818ff9_400007b7,
        64'hfe842703_f407dde3,
        64'hfe842783_fef42423,
        64'h87aa881f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783a4cd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_7ff000ef,
        64'hfb843503_90078593,
        64'h67ad863e_4681fe44,
        64'h2783fef4_22238fd9,
        64'h010007b7_fe442703,
        64'h00f71963_47a1873e,
        64'h4bdcfb84_378302f7,
        64'h10634789_873e0367,
        64'hc783fb84_3783fef4,
        64'h222340ff_87b7a689,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_05e010ef,
        64'hfb843503_70078593,
        64'h678d4601_4681a055,
        64'hfe042423_02e78aa3,
        64'h4709fb84_3783a031,
        64'h02e78aa3_4705fb84,
        64'h378300f7_08631aa0,
        64'h07930007_871bfe84,
        64'h2783fef4_242387aa,
        64'h94fff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_f3e52781,
        64'h8b892781_fe344783,
        64'hfef401a3_87aaa91f,
        64'hf0ef853e_02f00593,
        64'h43dcfb84_3783a821,
        64'hfef401a3_87aaaa9f,
        64'hf0ef853e_02f00593,
        64'h43dcfb84_3783af3f,
        64'hf0ef853e_02f00593,
        64'h460943dc_fb843783,
        64'h04f71863_47890007,
        64'h871bfec4_2783a129,
        64'hfef42623_478500f7,
        64'h06634789_0007871b,
        64'hfec42783_cf812781,
        64'hfec42783_fef42623,
        64'h87aa1340_10effb84,
        64'h35038007_85936785,
        64'h1aa00613_4681a189,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_15e010ef,
        64'hfb843503_45814601,
        64'h4681a19d_fef42623,
        64'h4785e789_27818ff9,
        64'h67c1fdc4_2703fcf4,
        64'h2e2387aa_a33ff0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfb84,
        64'h3783cb8d_47dcfb84,
        64'h378302f7_0e634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfb843783_a9754785,
        64'hc0e1ae23_4705f60f,
        64'hf0ef08a5_05130000,
        64'h451708a5_85930000,
        64'h45971620_0613a015,
        64'h04f71163_4789873e,
        64'h0367c783_fb843783,
        64'hcbd84711_fb843783,
        64'hc001ae23_a9f54785,
        64'hc0e1ae23_4705fa0f,
        64'hf0ef0ca5_05130000,
        64'h45170ca5_85930000,
        64'h45971610_0613a015,
        64'h04f71363_11178793,
        64'h111117b7_873e53dc,
        64'hfb843783_c001ae23,
        64'hcf91fb84_3783faa4,
        64'h3c230880_e0a2e486,
        64'h715d8082_61217442,
        64'h70e2853e_fec42783,
        64'hfe042623_be1ff0ef,
        64'h853e4591_20000613,
        64'h43dcfd84_3783c2e1,
        64'h9023474d_bf9ff0ef,
        64'h853e03a0_05934601,
        64'h43dcfd84_3783c0bf,
        64'hf0ef853e_03800593,
        64'h460143dc_fd843783,
        64'hc1dff0ef_853a0360,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c33f,
        64'hf0ef853a_03400593,
        64'heff78613_67c143d8,
        64'hfd843783_cc9ff0ef,
        64'h853e0280_05934641,
        64'h43dcfd84_3783cdbf,
        64'hf0ef853a_02900593,
        64'h863e0ff7_f7930017,
        64'he793feb4_478343d8,
        64'hfd843783_fe0405a3,
        64'ha019fef4_05a347a9,
        64'hc7892781_8ff90400,
        64'h07b7873e_579cfd84,
        64'h3783a005_fef405a3,
        64'h47b1c789_27818ff9,
        64'h020007b7_873e579c,
        64'hfd843783_a82dfef4,
        64'h05a347b9_c7892781,
        64'h8ff90100_07b7873e,
        64'h579cfd84_3783a8c5,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_0c0030ef,
        64'hfd843503_a8078593,
        64'h000627b7_b19ff0ef,
        64'h0c800513_00f71663,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cfd84_378302f7,
        64'h13634789_873e0367,
        64'hc783fd84_3783da3f,
        64'hf0ef853e_02900593,
        64'h463d43dc_fd843783,
        64'ha811db7f_f0ef853e,
        64'h02900593_463d43dc,
        64'hfd843783_00f71c63,
        64'h4789873e_0367c783,
        64'hfd843783_d798fd84,
        64'h37830007_871b87aa,
        64'hc8fff0ef_853e9381,
        64'h17822781_0407879b,
        64'h43dcfd84_378302e7,
        64'h8b23fd84_37830ff7,
        64'hf71387aa_d4fff0ef,
        64'h853e0fe0_059343dc,
        64'hfd843783_f3e52781,
        64'h8b852781_fea44783,
        64'hfef40523_87aadf1f,
        64'hf0ef853e_02f00593,
        64'h43dcfd84_3783a821,
        64'hfef40523_87aae09f,
        64'hf0ef853e_02f00593,
        64'h43dcfd84_3783e53f,
        64'hf0ef853e_02f00593,
        64'h460543dc_fd843783,
        64'hc0dff0ef_3e800513,
        64'he6dff0ef_853e0290,
        64'h05934601_43dcfd84,
        64'h3783a811_e81ff0ef,
        64'h853e0290_05934641,
        64'h43dcfd84_3783ac35,
        64'h4785c0e1_ae234705,
        64'ha33ff0ef_35c50513,
        64'h00004517_35c58593,
        64'h00004597_0b500613,
        64'ha01502f7_1e634789,
        64'h873e2781_0ff7f793,
        64'h278187aa_e0fff0ef,
        64'h853e0fe0_059343dc,
        64'hfd843783_0607b823,
        64'hfd843783_d7f84719,
        64'hfd843783_0607a223,
        64'hfd843783_02e78023,
        64'hfd843783_0207c703,
        64'hfd043783_cfd8fd84,
        64'h37834fd8_fd043783,
        64'hcf98fd84_37834f98,
        64'hfd043783_cbd8fd84,
        64'h37834bd8_fd043783,
        64'hcb98fd84_37834b98,
        64'hfd043783_c7d8fd84,
        64'h378347d8_fd043783,
        64'hd3d81117_071b1111,
        64'h1737fd84_3783c798,
        64'hfd843783_4798fd04,
        64'h3783c3d8_fcc42703,
        64'hfd843783_00e79023,
        64'hfd843783_0007d703,
        64'hfd043783_c001ae23,
        64'hae394785_c0e1ae23,
        64'h4705b15f_f0ef43e5,
        64'h05130000_451743e5,
        64'h85930000_45970b40,
        64'h0613a015_c3fdfd04,
        64'h3783c001_ae23c799,
        64'hfd843783_fcf42623,
        64'h87b2fcb4_3823fca4,
        64'h3c230080_f822fc06,
        64'h71398082_61056442,
        64'h60e20001_e8dff0ef,
        64'h853e85ba_fea44703,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_052387ba,
        64'hfef405a3_87b6fef4,
        64'h26238732_86ae87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h853e87aa_e7fff0ef,
        64'h853e9381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef405a3,
        64'h87bafef4_2623872e,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e20001_f39ff0ef,
        64'h853e85ba_fe845703,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_142387ba,
        64'hfef405a3_87b6fef4,
        64'h26238732_86ae87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h853e87aa_f1dff0ef,
        64'h853e9381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef405a3,
        64'h87bafef4_2623872e,
        64'h87aa1000_e822ec06,
        64'h11018082_61457422,
        64'h0001c398_fd442703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf42a23,
        64'h87aefca4_3c231800,
        64'hf4227179_80826145,
        64'h74220001_00e79023,
        64'hfd645703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf41b23_87aefca4,
        64'h3c231800_f4227179,
        64'h80826145_74220001,
        64'h00e78023_fd744703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf40ba3,
        64'h87aefca4_3c231800,
        64'hf4227179_80826105,
        64'h6462853e_2781439c,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61056462_853e93c1,
        64'h17c20007_d783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826105,
        64'h6462853e_0ff7f793,
        64'h0007c783_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61457422,
        64'h853efe84_3783fae7,
        64'hf5e34785_0007871b,
        64'hfe442783_fef42223,
        64'h2785fe44_2783a829,
        64'hfef43423_97ba0a67,
        64'h07131ffe_e717078a,
        64'h97ba078e_87bafe44,
        64'h670302f7_10632781,
        64'h2701fde4_57030007,
        64'hd78397ba_0d868713,
        64'h078a97ba_078e87ba,
        64'hfe446703_1ffee697,
        64'ha0b9fe04_2223fe04,
        64'h3423fcf4_1f2387aa,
        64'h1800f422_71798082,
        64'h61457402_70a20001,
        64'hfef768e3_fe043783,
        64'hfe843703_fea43423,
        64'hfbfff0ef_fef43023,
        64'h97bafe84_3783873e,
        64'h078a97ba_078a87ba,
        64'hfd843703_fea43423,
        64'hfdfff0ef_fca43c23,
        64'h1800f022_f4067179,
        64'h80820141_6422853e,
        64'h639c17e1_0200c7b7,
        64'h0800e422_11418082,
        64'h61096406_60a6853e,
        64'hfec42783_fef42623,
        64'h87aab38f_f0efc265,
        64'h0513ffff_f51785be,
        64'h567dfb84_3683fd04,
        64'h0793fe04_3703fcf4,
        64'h3c23fc04_3783fcf4,
        64'h3823fc84_3783fef4,
        64'h3023fd87_87930304,
        64'h07930314_34230304,
        64'h3023ec1c_e818e414,
        64'hfac43c23_fcb43023,
        64'hfca43423_0880e0a2,
        64'he4867119_80826145,
        64'h740270a2_853e87aa,
        64'hb9eff0ef_bf650513,
        64'hfffff517_fe843583,
        64'hfe043603_fd843683,
        64'hfd043703_fcd43823,
        64'hfcc43c23_feb43023,
        64'hfea43423_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_853e87aa,
        64'hbdeff0ef_c9450513,
        64'hfffff517_85be567d,
        64'hfd843683_fd043703,
        64'hfe840793_fcb43823,
        64'hfca43c23_1800f022,
        64'hf4067179_80826165,
        64'h744270e2_853efec4,
        64'h2783fef4_262387aa,
        64'hc1eff0ef_c7650513,
        64'hfffff517_fd843583,
        64'hfd043603_fc843683,
        64'h873efe04_3783fef4,
        64'h3023fd87_87930304,
        64'h07930314_34230304,
        64'h3023ec1c_e818e414,
        64'hfcc43423_fcb43823,
        64'hfca43c23_0080f822,
        64'hfc067159_80826125,
        64'h740270a2_853efec4,
        64'h2783fef4_262387aa,
        64'hc7eff0ef_cd650513,
        64'hfffff517_fd843583,
        64'h567dfd04_3683873e,
        64'hfe043783_fef43023,
        64'hfd078793_03040793,
        64'h03143423_03043023,
        64'hec1ce818_e414e010,
        64'hfcb43823_fca43c23,
        64'h1800f022_f406711d,
        64'h80826109_744270e2,
        64'h853efec4_2783fef4,
        64'h262387aa_cdaff0ef,
        64'hd9050513_fffff517,
        64'h85be567d_fc843683,
        64'hfd840793_fe043703,
        64'hfef43023_fc878793,
        64'h04040793_03143c23,
        64'h03043823_f41cf018,
        64'hec14e810_e40cfca4,
        64'h34230080_f822fc06,
        64'h71198082_610d644a,
        64'h60ea853e_2781fd84,
        64'h37839702_4501f904,
        64'h3583863e_f8843683,
        64'hf9843703_fd843783,
        64'ha01917fd_f8843783,
        64'h00f76663_f8843783,
        64'hfd843703_d8079963,
        64'h0007c783_f8043783,
        64'h0001f8f4_30230785,
        64'hf8043783_9702f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'h0007c503_f8043783,
        64'ha80df8f4_30230785,
        64'hf8043783_97020250,
        64'h0513f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_a8b9f8f4,
        64'h30230785_f8043783,
        64'hfca43c23_ba2ff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h87364781_484188ba,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442703,
        64'h86be639c_f6e43c23,
        64'h00878713_f7843783,
        64'ha089fca4_3c23cfcf,
        64'hf0eff984_3503f904,
        64'h3583fd84_3603f884,
        64'h36838736_47814841,
        64'h88bae03e_fe842783,
        64'he43efec4_2783fe44,
        64'h270386be_639cf6e4,
        64'h3c230087_8713f784,
        64'h3783c3b1_0ff7f793,
        64'hfbb44783_faf40da3,
        64'h4785fef4_26230217,
        64'he793fec4_2783fef4,
        64'h242347c1_a239f8f4,
        64'h30230785_f8043783,
        64'hfce7e7e3_2701fe84,
        64'h2703fce4_22230017,
        64'h871bfc44_27839702,
        64'h02000513_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_3783a00d,
        64'hcf8d2781_8b89fec4,
        64'h2783fbcd_fee42223,
        64'hfff7871b_fe442783,
        64'hd3e12781_4007f793,
        64'hfec42783_cf910007,
        64'hc783fc84_37839702,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h37830007_c503fce4,
        64'h34230017_8713fc84,
        64'h3783a03d_fce7e7e3,
        64'h2701fe84_2703fce4,
        64'h22230017_871bfc44,
        64'h27839702_02000513,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h3783a00d_e7a52781,
        64'h8b89fec4_2783fcf4,
        64'h222387b2_00d77363,
        64'h0006071b_0007869b,
        64'hfe442783_fc442603,
        64'hcf912781_4007f793,
        64'hfec42783_fcf42223,
        64'h87aa8aaf_f0effc84,
        64'h350385be_57fda011,
        64'hfe446783_c7812781,
        64'hfe442783_fcf43423,
        64'h639cf6e4_3c230087,
        64'h8713f784_3783a4a1,
        64'hf8f43023_0785f804,
        64'h3783fce7_e7e32701,
        64'hfe842703_fce42823,
        64'h0017871b_fd042783,
        64'h97020200_0513f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'ha00dcf8d_27818b89,
        64'hfec42783_9702f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'h0ff7f513_439cf6e4,
        64'h3c230087_8713f784,
        64'h3783fce7_e7e32701,
        64'hfe842703_fce42823,
        64'h0017871b_fd042783,
        64'h97020200_0513f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'ha00def8d_27818b89,
        64'hfec42783_fcf42823,
        64'h4785a631_f8f43023,
        64'h0785f804_3783fca4,
        64'h3c23e50f_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_36834781,
        64'h883688b2_e03efe84,
        64'h2783e43e_fec42783,
        64'hfe442603_fd446683,
        64'hfb446703_faf42a23,
        64'h2781439c_f6e43c23,
        64'h00878713_f7843783,
        64'ha8012781_93c117c2,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783cf81,
        64'h27810807_f793fec4,
        64'h2783a815_27810ff7,
        64'hf793439c_f6e43c23,
        64'h00878713_f7843783,
        64'hcf812781_0407f793,
        64'hfec42783_a841fca4,
        64'h3c23ee0f_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_36834781,
        64'h883688b2_e03efe84,
        64'h2783e43e_fec42783,
        64'hfe442603_fd446683,
        64'h6398f6e4_3c230087,
        64'h8713f784_3783c3b1,
        64'h27811007_f793fec4,
        64'h2783a8f9_fca43c23,
        64'h847ff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_47818836,
        64'h88b2e03e_fe842783,
        64'he43efec4_2783fe44,
        64'h2603fd44_66836398,
        64'hf6e43c23_00878713,
        64'hf7843783_c3b12781,
        64'h2007f793_fec42783,
        64'ha235fca4_3c23f7cf,
        64'hf0eff984_3503f904,
        64'h3583fd84_3603f884,
        64'h368387b6_883288ae,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442583,
        64'hfd446603_0ff7f693,
        64'h01f7d79b_fb042783,
        64'h93010207_97132781,
        64'h278140f7_07bb8f3d,
        64'hfb042703_41f7d79b,
        64'hfb042783_faf42823,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783a801,
        64'h27814107_d79b0107,
        64'h979b439c_f6e43c23,
        64'h00878713_f7843783,
        64'hcf912781_0807f793,
        64'hfec42783_a81d2781,
        64'h0ff7f793_439cf6e4,
        64'h3c230087_8713f784,
        64'h3783cf81_27810407,
        64'hf793fec4_2783a2cd,
        64'hfca43c23_833ff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h872e87ba_883688b2,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442603,
        64'hfd446683_0ff7f713,
        64'h93fdfa84_378385be,
        64'h8f998fb9_fa843783,
        64'h43f7d713_fa843783,
        64'hfaf43423_639cf6e4,
        64'h3c230087_8713f784,
        64'h3783c3bd_27811007,
        64'hf793fec4_2783ac89,
        64'hfca43c23_9bbff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h872e87ba_883688b2,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442603,
        64'hfd446683_0ff7f713,
        64'h93fdfa04_378385be,
        64'h8f998fb9_fa043783,
        64'h43f7d713_fa043783,
        64'hfaf43023_639cf6e4,
        64'h3c230087_8713f784,
        64'h3783c3bd_27812007,
        64'hf793fec4_278318f7,
        64'h1d630640_0793873e,
        64'h0007c783_f8043783,
        64'h00f70b63_06900793,
        64'h873e0007_c783f804,
        64'h3783fef4_26239bf9,
        64'hfec42783_c7912781,
        64'h4007f793_fec42783,
        64'hfef42623_9bcdfec4,
        64'h278300f7_07630640,
        64'h0793873e_0007c783,
        64'hf8043783_02f70063,
        64'h06900793_873e0007,
        64'hc783f804_3783fef4,
        64'h26230207_e793fec4,
        64'h278300f7_18630580,
        64'h0793873e_0007c783,
        64'hf8043783_fef42623,
        64'h9bbdfec4_2783fcf4,
        64'h2a2347a9_a809fcf4,
        64'h2a234789_00f71663,
        64'h06200793_873e0007,
        64'hc783f804_3783a035,
        64'hfcf42a23_47a100f7,
        64'h166306f0_0793873e,
        64'h0007c783_f8043783,
        64'ha099fcf4_2a2347c1,
        64'h00f71663_05800793,
        64'h873e0007_c783f804,
        64'h378300f7_0b630780,
        64'h0793873e_0007c783,
        64'hf8043783_878297ba,
        64'hee878793_00005797,
        64'h0007871b_439c97ba,
        64'hef878793_00005797,
        64'h00279713_93810206,
        64'h97936ce7_e3630530,
        64'h07930006_871bfdb7,
        64'h869b2781_0007c783,
        64'hf8043783_0001a011,
        64'h0001a021_0001a031,
        64'hf8f43023_0785f804,
        64'h3783fef4_26231007,
        64'he793fec4_2783a015,
        64'hf8f43023_0785f804,
        64'h3783fef4_26231007,
        64'he793fec4_2783a835,
        64'hf8f43023_0785f804,
        64'h3783fef4_26231007,
        64'he793fec4_2783a889,
        64'hf8f43023_0785f804,
        64'h3783fef4_26230407,
        64'he793fec4_278306f7,
        64'h16630680_0793873e,
        64'h0007c783_f8043783,
        64'hf8f43023_0785f804,
        64'h3783fef4_26230807,
        64'he793fec4_2783a079,
        64'hf8f43023_0785f804,
        64'h3783fef4_26232007,
        64'he793fec4_27830af7,
        64'h146306c0_0793873e,
        64'h0007c783_f8043783,
        64'hf8f43023_0785f804,
        64'h3783fef4_26231007,
        64'he793fec4_27838782,
        64'h97bafae7_87930000,
        64'h57970007_871b439c,
        64'h97bafbe7_87930000,
        64'h57970027_97139381,
        64'h02069793_0ee7e963,
        64'h47c90006_871bf987,
        64'h869b2781_0007c783,
        64'hf8043783_f8f43023,
        64'h0785f804_3783fef4,
        64'h22232781_47810007,
        64'h53630007_871bfbc4,
        64'h2783faf4_2e23439c,
        64'hf6e43c23_00878713,
        64'hf7843783_02f71a63,
        64'h02a00793_873e0007,
        64'hc783f804_3783a091,
        64'hfef42223_87aaf86f,
        64'hf0ef853e_f8040793,
        64'hcb9187aa_f54ff0ef,
        64'h853e0007_c783f804,
        64'h3783f8f4_30230785,
        64'hf8043783_fef42623,
        64'h4007e793_fec42783,
        64'h08f71063_02e00793,
        64'h873e0007_c783f804,
        64'h3783fe04_2223f8f4,
        64'h30230785_f8043783,
        64'hfef42423_fc042783,
        64'ha029fef4_24232781,
        64'h40f007bb_fc042783,
        64'hfef42623_0027e793,
        64'hfec42783_0207d063,
        64'h2781fc04_2783fcf4,
        64'h2023439c_f6e43c23,
        64'h00878713_f7843783,
        64'h04f71763_02a00793,
        64'h873e0007_c783f804,
        64'h3783a8b9_fef42423,
        64'h87aa833f_f0ef853e,
        64'hf8040793_cb9187aa,
        64'h801ff0ef_853e0007,
        64'hc783f804_3783fe04,
        64'h2423f385_2781fe04,
        64'h27830001_fe042023,
        64'ha021fef4_20234785,
        64'hf8f43023_0785f804,
        64'h3783fef4_26230107,
        64'he793fec4_2783a01d,
        64'hfef42023_4785f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0087e793,
        64'hfec42783_a091fef4,
        64'h20234785_f8f43023,
        64'h0785f804_3783fef4,
        64'h26230047_e793fec4,
        64'h2783a08d_fef42023,
        64'h4785f8f4_30230785,
        64'hf8043783_fef42623,
        64'h0027e793_fec42783,
        64'ha041fef4_20234785,
        64'hf8f43023_0785f804,
        64'h3783fef4_26230017,
        64'he793fec4_27838782,
        64'h97ba1627_87930000,
        64'h57970007_871b439c,
        64'h97ba1727_87930000,
        64'h57970027_97139381,
        64'h02069793_0ce7e063,
        64'h47c10006_871bfe07,
        64'h869b2781_0007c783,
        64'hf8043783_fe042623,
        64'hf8f43023_0785f804,
        64'h37832270_006ff8f4,
        64'h30230785_f8043783,
        64'h9702f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_0007c503,
        64'hf8043783_02f70b63,
        64'h02500793_873e0007,
        64'hc783f804_378326b0,
        64'h006ff8f4_3c238667,
        64'h87930000_07972607,
        64'h9de3f904_3783fc04,
        64'h3c23f6e4_3c23f8d4,
        64'h3023f8c4_3423f8b4,
        64'h3823f8a4_3c231100,
        64'he922ed06_71358082,
        64'h610d644a_60ea853e,
        64'h87aab47f_f0effb84,
        64'h3503fb04_3583fa84,
        64'h3603fa04_3683fe84,
        64'h37838836_88b2e03e,
        64'hf9042783_e43e401c,
        64'he83e441c_fc040713,
        64'hf9744683_0007861b,
        64'hf8843783_f6e7ffe3,
        64'h47fdfe84_3703c791,
        64'hf9843783_f8f43c23,
        64'h02f757b3_f8843783,
        64'hf9843703_fcf70823,
        64'h9736ff04_0693fed4,
        64'h34230017_0693fe84,
        64'h37030ff7_f79337d9,
        64'h0ff7f793_9fb9fe74,
        64'h47030610_0793a019,
        64'h04100793_c7812781,
        64'h0207f793_441ca01d,
        64'h0ff7f793_0307879b,
        64'hfe744783_00e7e963,
        64'h47a50ff7_f713fe74,
        64'h4783fef4_03a302f7,
        64'h77b3f884_3783f984,
        64'h3703c7c1_f9843783,
        64'hc7812781_4007f793,
        64'h441cc41c_9bbd441c,
        64'he781f984_3783fe04,
        64'h3423f8f4_282387ba,
        64'hf8f40ba3_8746f904,
        64'h3423f8e4_3c23fad4,
        64'h3023fac4_3423fab4,
        64'h3823faa4_3c231100,
        64'he922ed06_71358082,
        64'h610d644a_60ea853e,
        64'h87aac5ff_f0effb84,
        64'h3503fb04_3583fa84,
        64'h3603fa04_3683fe84,
        64'h37838836_88b2e03e,
        64'hf9042783_e43e401c,
        64'he83e441c_fc040713,
        64'hf9744683_0007861b,
        64'hf8843783_f6e7ffe3,
        64'h47fdfe84_3703c791,
        64'hf9843783_f8f43c23,
        64'h02f757b3_f8843783,
        64'hf9843703_fcf70823,
        64'h9736ff04_0693fed4,
        64'h34230017_0693fe84,
        64'h37030ff7_f79337d9,
        64'h0ff7f793_9fb9fe74,
        64'h47030610_0793a019,
        64'h04100793_c7812781,
        64'h0207f793_441ca01d,
        64'h0ff7f793_0307879b,
        64'hfe744783_00e7e963,
        64'h47a50ff7_f713fe74,
        64'h4783fef4_03a302f7,
        64'h77b3f884_3783f984,
        64'h3703c7c1_f9843783,
        64'hc7812781_4007f793,
        64'h441cc41c_9bbd441c,
        64'he781f984_3783fe04,
        64'h3423f8f4_282387ba,
        64'hf8f40ba3_8746f904,
        64'h3423f8e4_3c23fad4,
        64'h3023fac4_3423fab4,
        64'h3823faa4_3c231100,
        64'he922ed06_71358082,
        64'h61616406_60a6853e,
        64'h87aac65f_f0effe84,
        64'h3503fe04_3583fd84,
        64'h3603fd04_3683fc84,
        64'h3703fc04_3783883e,
        64'h88ba441c_481800e7,
        64'h80230200_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'hcf912781_8ba1481c,
        64'ha01500e7_802302b0,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_cf992781,
        64'h8b91481c_a0a100e7,
        64'h802302d0_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'hcf990ff7_f793fbf4,
        64'h478306e7_e86347fd,
        64'hfc043703_00e78023,
        64'h03000713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_378300e7,
        64'hef6347fd_fc043703,
        64'h00e78023_06200713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h378300e7_ef6347fd,
        64'hfc043703_02f71463,
        64'h47890007_871bfb84,
        64'h2783a815_00e78023,
        64'h05800713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_378302e7,
        64'he06347fd_fc043703,
        64'hc7852781_0207f793,
        64'h481c02f7_1a6347c1,
        64'h0007871b_fb842783,
        64'ha88d00e7_80230780,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_02e7e063,
        64'h47fdfc04_3703e785,
        64'h27810207_f793481c,
        64'h02f71a63_47c10007,
        64'h871bfb84_2783fcf4,
        64'h302317fd_fc043783,
        64'h00f71763_47c10007,
        64'h871bfb84_2783cf89,
        64'hfc043783_fcf43023,
        64'h17fdfc04_378302f7,
        64'h1663fc04_37030084,
        64'h678300f7_0863fc04,
        64'h37030004_6783c3a9,
        64'hfc043783_e7a12781,
        64'h4007f793_481c1207,
        64'h83632781_8bc1481c,
        64'hfce7f6e3_47fdfc04,
        64'h370300f7_7763fc04,
        64'h37030084_6783cf81,
        64'h27818b85_481c00e7,
        64'h80230300_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'ha831fce7_fae347fd,
        64'hfc043703_02f77563,
        64'hfc043703_00046783,
        64'h00e78023_03000713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h3783a831_c41c37fd,
        64'h441cc395_27818bb1,
        64'h481ce789_0ff7f793,
        64'hfbf44783_cb9d2781,
        64'h8b85481c_cf9d2781,
        64'h441cebd1_27818b89,
        64'h481cfaf4_2c2387ba,
        64'hfaf40fa3_874687c2,
        64'hfcf43023_fce43423,
        64'hfcd43823_fcc43c23,
        64'hfeb43023_fea43423,
        64'h0880e0a2_e486715d,
        64'h80826125_644660e6,
        64'h853efc84_3783fcf7,
        64'h69e3fac4_67838f1d,
        64'hfe043783_fc843703,
        64'h97020200_0513fd04,
        64'h3583863e_fc043683,
        64'hfd843703_fce43423,
        64'h00178713_fc843783,
        64'ha00dcb9d_27818b89,
        64'hfa842783_f7e1fb04,
        64'h37839702_fd043583,
        64'h863efc04_3683fd84,
        64'h3703fce4_34230017,
        64'h8713fc84_37830007,
        64'hc50397ba_fb043783,
        64'hfb843703_faf43823,
        64'h17fdfb04_3783a81d,
        64'hfcf767e3_fe843703,
        64'hfac46783_fef43423,
        64'h0785fe84_37839702,
        64'h02000513_fd043583,
        64'h863efc04_3683fd84,
        64'h3703fce4_34230017,
        64'h8713fc84_3783a035,
        64'hfef43423_fb043783,
        64'hefa52781_8b85fa84,
        64'h2783e3c9_27818b89,
        64'hfa842783_fef43023,
        64'hfc843783_faf42423,
        64'h87bafaf4_26238746,
        64'h87c2faf4_3823fae4,
        64'h3c23fcd4_3023fcc4,
        64'h3423fcb4_3823fca4,
        64'h3c231080_e8a2ec86,
        64'h711d8082_61457402,
        64'h70a2853e_fec42783,
        64'hffc587aa_f6dff0ef,
        64'h853e0007_c783639c,
        64'hfd843783_fef42623,
        64'hfd07879b_27819fb9,
        64'h27810007_c783e290,
        64'hfd843683_00178613,
        64'h639cfd84_37830007,
        64'h871b0017_979b9fb9,
        64'h0027979b_87bafec4,
        64'h2703a825_fe042623,
        64'hfca43c23_1800f022,
        64'hf4067179_80826105,
        64'h6462853e_0ff7f793,
        64'h8b854781_a0114785,
        64'h00e7e463_03900793,
        64'h0ff7f713_fef44783,
        64'h00e7fc63_02f00793,
        64'h0ff7f713_fef44783,
        64'hfef407a3_87aa1000,
        64'hec221101_80826145,
        64'h7422853e_278140f7,
        64'h07b3fd84_3783fe84,
        64'h3703f3e5_fce43823,
        64'hfff78713_fd043783,
        64'hcb810007_c783fe84,
        64'h3783fef4_34230785,
        64'hfe843783_a031fef4,
        64'h3423fd84_3783fcb4,
        64'h3823fca4_3c231800,
        64'hf4227179_80826145,
        64'h740270a2_00019682,
        64'h853e85ba_fef44783,
        64'h6798fe04_37836394,
        64'hfe043783_cf810ff7,
        64'hf793fef4_4783fef4,
        64'h07a3fcd4_3823fcc4,
        64'h3c23feb4_302387aa,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h00018e7f_f0ef853e,
        64'hfef44783_c7910ff7,
        64'hf793fef4_4783fef4,
        64'h07a3fcd4_3823fcc4,
        64'h3c23feb4_302387aa,
        64'h1800f022_f4067179,
        64'h80826145_74220001,
        64'hfef407a3_fcd43823,
        64'hfcc43c23_feb43023,
        64'h87aa1800_f4227179,
        64'h80826145_74220001,
        64'h00e78023_fef44703,
        64'h97bafd84_3783fe04,
        64'h370300f7_7b63fd04,
        64'h3783fd84_3703fef4,
        64'h07a3fcd4_3823fcc4,
        64'h3c23feb4_302387aa,
        64'h1800f422_71798082,
        64'h610d690a_64aa644a,
        64'h60eaf604_0113853e,
        64'h8126814a_47812b00,
        64'h10ef9ea5_05130000,
        64'h6517a801_57f92c00,
        64'h10ef7aa5_05130000,
        64'h551785be_fac42783,
        64'h2d2010ef_7a450513,
        64'h00005517_c3952781,
        64'hfac42783_faf42623,
        64'h87aab63f_f0eff684,
        64'h350385be_863af644,
        64'h27032781_739cf804,
        64'h37833040_10efa265,
        64'h05130000_6517f8f4,
        64'h3023f884_3783eae7,
        64'hd2e3478d_0007871b,
        64'hfd042783_fcf42823,
        64'h2785fd04_27833300,
        64'h10ef8725_05130000,
        64'h6517fce7_d6e30470,
        64'h07930007_871bfdc4,
        64'h2783fcf4_2e232785,
        64'hfdc42783_356010ef,
        64'h9f050513_00006517,
        64'h85be2781_0387c783,
        64'h97bafdc4_2783f784,
        64'h3703a02d_fc042e23,
        64'h37a010ef_a8450513,
        64'h00006517_386010ef,
        64'ha7850513_00006517,
        64'h85be7b9c_f7843783,
        64'h39a010ef_a7450513,
        64'h00006517_85be779c,
        64'hf7843783_3ae010ef,
        64'ha7050513_00006517,
        64'h85be739c_f7843783,
        64'hfce7d7e3_47bd0007,
        64'h871bfd84_2783fcf4,
        64'h2c232785_fd842783,
        64'h3da010ef_a7450513,
        64'h00006517_85be2781,
        64'h0107c783_97bafd84,
        64'h2783f784_3703a02d,
        64'hfc042c23_3fe010ef,
        64'haa050513_00006517,
        64'hfce7d7e3_47bd0007,
        64'h871bfd44_2783fcf4,
        64'h2a232785_fd442783,
        64'h422010ef_abc50513,
        64'h00006517_85be2781,
        64'h0007c783_97bafd44,
        64'h2783f784_3703a02d,
        64'hfc042a23_446010ef,
        64'hac050513_00006517,
        64'h452010ef_ab450513,
        64'h00006517_85befd04,
        64'h2783f6f4_3c2397ba,
        64'h27010077_171bfd04,
        64'h2703f884_3783aa91,
        64'hfc042823_aac957f9,
        64'h482010ef_ac450513,
        64'h00006517_85befac4,
        64'h27834940_10ef9665,
        64'h05130000_6517c395,
        64'h2781fac4_2783faf4,
        64'h262387aa_d25ff0ef,
        64'h853a85be_46052781,
        64'h67bcfa04_3783f884,
        64'h3703f8f4_34230007,
        64'h8793878a_40f10133,
        64'h07928391_07bdf8e4,
        64'h3823177d_873e893a,
        64'h870afc04_37834e80,
        64'h10efb0a5_05130000,
        64'h651785be_4bfcfa04,
        64'h37834fc0_10efafe5,
        64'h05130000_651785be,
        64'h4bbcfa04_37835100,
        64'h10efaea5_05130000,
        64'h651785be_67bcfa04,
        64'h37835240_10efae65,
        64'h05130000_651785be,
        64'h739cfa04_37835380,
        64'h10efae25_05130000,
        64'h651785be_6f9cfa04,
        64'h378354c0_10efade5,
        64'h05130000_651785be,
        64'h4bdcfa04_37835600,
        64'h10efada5_05130000,
        64'h651785be_4b9cfa04,
        64'h37835740_10efad65,
        64'h05130000_651785be,
        64'h47dcfa04_37835880,
        64'h10efad25_05130000,
        64'h651785be_479cfa04,
        64'h378359c0_10efade5,
        64'h05130000_6517fce7,
        64'hd7e3479d_0007871b,
        64'hfcc42783_fcf42623,
        64'h2785fcc4_27835c00,
        64'h10efafa5_05130000,
        64'h651785be_27810007,
        64'hc78397ba_f9843703,
        64'hfcc42783_a02dfc04,
        64'h2623f8f4_3c23fa04,
        64'h37835ec0_10efb165,
        64'h05130000_65175f80,
        64'h10efb025_05130000,
        64'h6517faf4_3023fb04,
        64'h3783a68d_57f96100,
        64'h10efafa5_05130000,
        64'h651785be_fac42783,
        64'h622010ef_af450513,
        64'h00006517_c3952781,
        64'hfac42783_faf42623,
        64'h87aaeb3f_f0ef853e,
        64'h45854605_fb043783,
        64'hfaf43823_00078793,
        64'h878a40f1_01330792,
        64'h839107bd_fae43c23,
        64'h177d873e_fc043783,
        64'hfcf43023_20000793,
        64'h672010ef_b2c50513,
        64'h00006517_aed157fd,
        64'h682010ef_b1450513,
        64'h00006517_cb892781,
        64'hfc842783_fcf42423,
        64'h87aae5bf_f0ef84be,
        64'h878af6f4_222387ae,
        64'hf6a43423_1100e14a,
        64'he526e922_ed067135,
        64'h80826145_740270a2,
        64'h853e4781_a01157fd,
        64'h6ca010ef_b3c50513,
        64'h00006517_85befe44,
        64'h2783cf81_2781fe44,
        64'h2783fef4_222387aa,
        64'h760030ef_26450513,
        64'h1fff0517_85be863a,
        64'hfe843683_fd442783,
        64'hfd042703_fae7e0e3,
        64'h678d0007_871bfd04,
        64'h2783fef4_342397ba,
        64'h006007b7_fe843703,
        64'hfcf42823_9fb977f5,
        64'hfd042703_a0b557fd,
        64'h732010ef_ba450513,
        64'h00006517_85befe04,
        64'h2783cf81_2781fe04,
        64'h2783fef4_202387aa,
        64'h7c8030ef_2cc50513,
        64'h1fff0517_85be660d,
        64'hfe843683_fd442783,
        64'ha8a1fef4_3423fd84,
        64'h3783fcf4_282387ba,
        64'hfcf42a23_873287ae,
        64'hfca43c23_1800f022,
        64'hf4067179_80826105,
        64'h644260e2_853e4781,
        64'h79a010ef_bec50513,
        64'h00006517_a80157f5,
        64'h7aa010ef_bcc50513,
        64'h00006517_85befe44,
        64'h2783cf81_2781fe44,
        64'h2783fef4_222387aa,
        64'h53c020ef_34450513,
        64'h1fff0517_a08157f9,
        64'h7da010ef_bd450513,
        64'h00006517_85befe44,
        64'h2783cf81_2781fe44,
        64'h2783fef4_222387aa,
        64'h4ab010ef_37450513,
        64'h1fff0517_fe843583,
        64'h863e43dc_fe843783,
        64'ha8b557fd_017010ef,
        64'hbf050513_00006517,
        64'heb89fe84_3783fea4,
        64'h34232890_10ef4501,
        64'h033010ef_bf450513,
        64'h00006517_1000e822,
        64'hec061101_80826145,
        64'h740270a2_0001eb9f,
        64'hf0ef0107_851307fa,
        64'h478d0200_0593ec9f,
        64'hf0ef0087_851307fa,
        64'h478d0c70_0593ed9f,
        64'hf0ef00c7_851307fa,
        64'h478d458d_ee7ff0ef,
        64'h00478513_07fa478d,
        64'h85be0ff7_f7932781,
        64'h0087d79b_fec42783,
        64'hf03ff0ef_01e79513,
        64'h478d85be_0ff7f793,
        64'hfec42783_f17ff0ef,
        64'h00c78513_07fa478d,
        64'h08000593_f27ff0ef,
        64'h00478513_07fa478d,
        64'h4581fef4_262302f7,
        64'h57bbfdc4_27032781,
        64'h0047979b_fd842783,
        64'hfcf42c23_87bafcf4,
        64'h2e23872e_87aa1800,
        64'hf022f406_71798082,
        64'h61056442_60e20001,
        64'hf6bff0ef_01e79513,
        64'h478d85be_fef44783,
        64'hdfed87aa_fc9ff0ef,
        64'h0001fef4_07a387aa,
        64'h1000e822_ec061101,
        64'h80820141_640260a2,
        64'h853e2781_0207f793,
        64'h278187aa_fd3ff0ef,
        64'h01478513_07fa478d,
        64'h0800e022_e4061141,
        64'h80826105_6462853e,
        64'h0ff7f793_0007c783,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61457422_000100e7,
        64'h8023fd74_4703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_0ba387ae,
        64'hfca43c23_1800f422,
        64'h7179a001_19f010ef,
        64'hd3850513_00006517,
        64'h84023025_85930000,
        64'h65971000_0437eb81,
        64'h2781fe44_27831c10,
        64'h10efd325_05130000,
        64'h6517fce7_d7e347bd,
        64'h0007871b_fe842783,
        64'hfef42423_2785fe84,
        64'h27831e50_10efd765,
        64'h05130000_651785be,
        64'h27810007_c78397ba,
        64'hfd843703_fe842783,
        64'ha02dfe04_24232090,
        64'h10efd825_05130000,
        64'h65171000_05b7fcf4,
        64'h3c231000_07b7fef4,
        64'h222387aa_370000ef,
        64'h10000537_65a12310,
        64'h10efda25_05130000,
        64'h6517fae7_d0e34789,
        64'h0007871b_fec42783,
        64'hfef42623_2785fec4,
        64'h27832550_10efdbe5,
        64'h05130000_651785b6,
        64'h863e43dc_97ba078e,
        64'hda470713_fec42783,
        64'h1fff0717_439497ba,
        64'hdb678793_070efec4,
        64'h27031fff_07972890,
        64'h10efdea5_05130000,
        64'h65174a70_10ef2407,
        64'h8513000f_47b7a8a1,
        64'hfe042623_2a7010ef,
        64'hde050513_00006517,
        64'h1be000ef_a0078513,
        64'h026267b7_20078593,
        64'h67f11800_f022f406,
        64'h7179f67f_f06f0141,
        64'h60a2e0a0_80e7ffff,
        64'h0097e406_7b850513,
        64'h80858593_11412000,
        64'h05372000_15b7c38d,
        64'h00078793_000007b7,
        64'h80828082_01416402,
        64'h60a280f4_00234785,
        64'he40080e7_ffff0097,
        64'h7b850513_20000537,
        64'hcb890007_87930000,
        64'h07b7f97f_f0ef843e,
        64'he406e022_1141eb1d,
        64'h8007c703_200017b7,
        64'h80828302_7b850513,
        64'h00030563_00030313,
        64'h00000337_c99102f5,
        64'hc5b34789_858d8d9d,
        64'h7b850793_7b878593,
        64'h20000537_200007b7,
        64'h80828302_7b850513,
        64'h00030563_00030313,
        64'h00000337_00e78b63,
        64'h7b878793_7b850713,
        64'h200007b7_20000537,
        64'h80823b50_506f0d00,
        64'h00ef4601_002c4502,
        64'h42d050ef_3bb050ef,
        64'hbf050513_00006517,
        64'h49f050ef_45818e09,
        64'hef060613_3fff0617,
        64'h6b050513_1fff0517,
        64'hea818193_1fff1197,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00048067,
        64'h100004b7_54c58593,
        64'h00006597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h192000ef_f9410113,
        64'h3fff0117_4f1050ef,
        64'hfeb56ce3_00450513,
        64'h00052023_00b57863,
        64'hc2218593_76c50513,
        64'h1fff0517_fec5e8e3,
        64'h00458593_00450513,
        64'h0055a023_00052283,
        64'h00c5fc63_78c60613,
        64'h1fff0617_fdc58593,
        64'h1fff0597_1e450513,
        64'h00007517_f9418193,
        64'h1fff1197_09249263,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
