/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 3134;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00000058_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000058_36313025,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000058_36313025,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_58323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h000a5838_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h000a5838_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_0000000a,
        64'h58363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h0000000a_58363130,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h0000000a_58363130,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_0a583830,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_0a583830,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_0a583830,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_0a583830,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h0000000a_58363130,
        64'h25202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h00000000_0a642520,
        64'h3a737574_61747320,
        64'h2c64656c_69616620,
        64'h64616552_20304453,
        64'h00000000_0a216465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a6425,
        64'h203a7375_74617473,
        64'h202c6465_6c696166,
        64'h206e6f69_74617a69,
        64'h6c616974_696e6920,
        64'h64726163_20304453,
        64'h0000000a_6425203a,
        64'h73757461_7473202c,
        64'h64656c69_6166206c,
        64'h61697469_6e692067,
        64'h69666e6f_63204453,
        64'h00000000_0000000a,
        64'h2164656c_69616620,
        64'h6769666e_6f632070,
        64'h756b6f6f_6c204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000a2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd0080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h08090000_38000000,
        64'hda0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000a001,
        64'h80cfc0ef_1c450513,
        64'h00001517_84025be5,
        64'h85930000_05971000,
        64'h0437e901_da6fb0ef,
        64'h10000537_65a1f475,
        64'h834fc0ef_347d1e65,
        64'h05130000_1517930f,
        64'hc0ef8526_24048493,
        64'h442984ef_c0ef000f,
        64'h44b71da5_05130000,
        64'h1517cecf_b0efe426,
        64'he822ec06_a0050513,
        64'h20058593_11010262,
        64'h653765f1_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623978f,
        64'hc0ef4505_a031fef4,
        64'h26234785_e7892781,
        64'h0807f793_278187aa,
        64'ha31fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'h0001a011_f6e7fee3,
        64'h02700793_0ff7f713,
        64'hfe944783_fef404a3,
        64'h2785fe94_4783cf99,
        64'h27810407_f7932781,
        64'h87aaa6bf_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h3783a0ad_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'ha61fd0ef_fd843503,
        64'h50078593_67854601,
        64'h4685a829_fef42623,
        64'h87aaa7bf_d0effd84,
        64'h35033007_85936785,
        64'h46014685_00f71f63,
        64'h4785873e_0347c783,
        64'hfd843783_a8adfe04,
        64'h04a3a34f_c0ef4505,
        64'hb13fe0ef_853e03e0,
        64'h0593863a_fe645703,
        64'h43dcfd84_3783fef4,
        64'h13230407_e793fe64,
        64'h5783fef4_132387aa,
        64'hb01fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'h66e79923_47410000,
        64'h0797b55f_e0ef853e,
        64'h4591863a_fea45703,
        64'h43dcfd84_3783fef4,
        64'h15238ff9_17fd6785,
        64'hfea45703_fef41523,
        64'h0017979b_fea45783,
        64'haa354785_6ae7a523,
        64'h47050000_07979caf,
        64'hc0ef75a5_05130000,
        64'h05177525_85930000,
        64'h059748e0_0613a025,
        64'h02f71c63_478d873e,
        64'h0377c783_fd843783,
        64'hfef41523_04000793,
        64'h6e07a223_00000797,
        64'ha2514785_6ee7a923,
        64'h47050000_0797a12f,
        64'hc0ef7a25_05130000,
        64'h051779a5_85930000,
        64'h059748d0_0613a025,
        64'h04f71763_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_7207a423,
        64'h00000797_c385fd84,
        64'h3783fca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'hb8ffe0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_c4ffe0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe842783,
        64'ha83dfef4_26234785,
        64'hc73fe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe84,
        64'h2703fef4_242387aa,
        64'hc61fe0ef_853e0300,
        64'h059343dc_fd843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aac57f,
        64'hd0effd84_35036000,
        64'h0593863e_4681fd44,
        64'h2783fcf4_2a2387ae,
        64'hfca43c23_1800f022,
        64'hf4067179_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aac55f,
        64'he0ef853e_93811782,
        64'h278127c1_43dcfc84,
        64'h3783d15f_e0ef853e,
        64'h03000593_460943dc,
        64'hfc843783_dfc52781,
        64'h8b89fdc4_2783a83d,
        64'hfef42623_4785d39f,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfc843783_c3852781,
        64'h8ff967a1_fdc42703,
        64'hfcf42e23_87aad27f,
        64'he0ef853e_03000593,
        64'h43dcfc84_3783a8bd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_d1dfd0ef,
        64'hfc843503_80078593,
        64'h6785863e_4685fe44,
        64'h27838ce7_92234745,
        64'h00001797_f56fe0ef,
        64'hfc843503_85befc04,
        64'h36032781_fe245783,
        64'hdbbfe0ef_853e4591,
        64'h863afe04_570343dc,
        64'hfc843783_fef41023,
        64'h8ff917fd_6785fe04,
        64'h5703fef4_10232000,
        64'h0793fef4_11234785,
        64'hfce7dee3_1ff00793,
        64'h0007871b_fe842783,
        64'hfef42423_2785fe84,
        64'h27830007_802397ba,
        64'hfc043703_fe842783,
        64'ha2154785_92e7ad23,
        64'h47050000_1797c5af,
        64'hc0ef9ea5_05130000,
        64'h15179e25_85930000,
        64'h159735d0_0613a081,
        64'hfe042423_9607a023,
        64'h00001797_aaa14785,
        64'h96e7a723_47050000,
        64'h1797c8ef_c0efa1e5,
        64'h05130000_1517a165,
        64'h85930000_159735c0,
        64'h0613a025_02f71d63,
        64'h11178793_111117b7,
        64'h873e53dc_fc843783,
        64'h9a07a223_00001797,
        64'hc385fc84_3783fe04,
        64'h2223fcb4_3023fca4,
        64'h34230080_f822fc06,
        64'h71398082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_a019fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aae63f_d0effd84,
        64'h3503a007_859367ad,
        64'h46014681_a03dfef4,
        64'h26234785_a82d4785,
        64'ha0e7a723_47050000,
        64'h1797d2ef_c0efabe5,
        64'h05130000_1517ab65,
        64'h85930000_159732d0,
        64'h0613a025_cb8d2781,
        64'hfec42783_fef42623,
        64'h87aaeb3f_d0effd84,
        64'h35037007_8593678d,
        64'h863e4681_4bbcfd84,
        64'h3783a407_ab230000,
        64'h1797a841_4785a6e7,
        64'ha2234705_00001797,
        64'hd84fc0ef_b1450513,
        64'h00001517_b0c58593,
        64'h00001597_32c00613,
        64'ha02504f7_1e631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783a807,
        64'had230000_1797c385,
        64'hfd843783_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efe84_2783fe04,
        64'h2423fa5f_e0ef853a,
        64'h02c00593_863e93c1,
        64'h17c20047_e793fe44,
        64'h578343d8_fd843783,
        64'hfef41223_87aaf8ff,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783d3e5,
        64'h27818b89_2781fe64,
        64'h5783fef4_132387aa,
        64'hfb1fe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'ha821fef4_132387aa,
        64'hfc9fe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'h812ff0ef_853e02c0,
        64'h0593863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12230017_e79393c1,
        64'h17c28fd9_fe445783,
        64'hfec45703_fef41623,
        64'hf007f793_fec45783,
        64'hfef41623_0087979b,
        64'hfec45783_fef41223,
        64'h0ff7f793_fe445783,
        64'hfef41223_87aa82ef,
        64'hf0ef853e_02c00593,
        64'h43dcfd84_3783a0a5,
        64'h87aff0ef_853e02c0,
        64'h0593863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12230017_e79393c1,
        64'h17c28fd9_fe445783,
        64'h93410307_97138fd9,
        64'hfe245783_fec45703,
        64'hfef41623_f007f793,
        64'hfec45783_fef41623,
        64'h0087979b_fec45783,
        64'hfef41123_0c07f793,
        64'hfe245783_fef41123,
        64'h0067979b_fe245783,
        64'hfef41123_0087d79b,
        64'hfec45783_fef41223,
        64'h03f7f793_fe445783,
        64'hfef41223_87aa8c6f,
        64'hf0ef853e_02c00593,
        64'h43dcfd84_378308f7,
        64'h1e634789_873e0367,
        64'hc783fd84_3783a249,
        64'hfef42423_478500e7,
        64'hf6631000_07930007,
        64'h871bfee4_5783fae7,
        64'hfee31000_07930007,
        64'h871bfee4_5783fef4,
        64'h17230017_979bfee4,
        64'h5783a839_fef41623,
        64'h0017d79b_fee45783,
        64'h00e7e963_2781fd44,
        64'h27830007_871b02f7,
        64'h57bb2781_fee45783,
        64'h4798fd84_3783a82d,
        64'hfef41723_4785a2ed,
        64'hfef42423_478506e7,
        64'hfa637fe0_07930007,
        64'h871bfee4_5783fae7,
        64'hffe37fe0_07930007,
        64'h871bfee4_5783fef4,
        64'h17232785_fee45783,
        64'ha831fef4_16230017,
        64'hd79bfee4_578300e7,
        64'he9632781_fd442783,
        64'h0007871b_02f757bb,
        64'h2781fee4_57834798,
        64'hfd843783_a825fef4,
        64'h17234785_ac914785,
        64'hd0e7ab23_47050000,
        64'h1797837f_c0efdc65,
        64'h05130000_1517dbe5,
        64'h85930000_15972b80,
        64'h0613a025_08f71963,
        64'h4789873e_0367c783,
        64'hfd843783_a26ff0ef,
        64'h853e02c0_0593863a,
        64'hfe445703_43dcfd84,
        64'h3783fef4_12239be9,
        64'hfe445783_fef41223,
        64'h87aaa12f_f0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783d607_af230000,
        64'h1797a4e9_4785d8e7,
        64'ha6234705_00001797,
        64'h8adfc0ef_e3c50513,
        64'h00001517_e3458593,
        64'h00001597_2b700613,
        64'ha02506f7_1e631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783dc07,
        64'ha1230000_1797c385,
        64'hfd843783_fe041623,
        64'hfcf42a23_87aefca4,
        64'h3c231800_f022f406,
        64'h71798082_61657406,
        64'h70a6853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_a32ff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_f9843783,
        64'hb72ff0ef_853e0280,
        64'h0593863a_0ff77713,
        64'hfe442703_43dcf984,
        64'h3783fef4_22230047,
        64'he793fe44_2783fef4,
        64'h222387aa_b64ff0ef,
        64'h853e0280_059343dc,
        64'hf9843783_a57fc0ef,
        64'h3e800513_a09dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa7300_00eff984,
        64'h350302f7_1163479d,
        64'h873e57fc_f9843783,
        64'ha849fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa0b80,
        64'h00eff984_350385be,
        64'h5f9cf984_3783b88f,
        64'hf0ef853e_03000593,
        64'h460943dc_f9843783,
        64'hdfc52781_8b89fe44,
        64'h2783a8d1_fef42623,
        64'h4785bacf_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_f9843783,
        64'hc3852781_8ff967a1,
        64'hfe442703_fef42223,
        64'h87aab9af_f0ef853e,
        64'h03000593_43dcf984,
        64'h3783aa11_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hb90fe0ef_f9843503,
        64'h60000593_863e4681,
        64'hfe842783_df985007,
        64'h071b0319_7737f984,
        64'h3783fef4_24231007,
        64'h879b03b9_07b7a831,
        64'hdf985007_071b0319,
        64'h7737f984_3783fef4,
        64'h24231007_879b03b9,
        64'h07b702f7_10634791,
        64'h873e57fc_f9843783,
        64'ha099df98_2007071b,
        64'h0bebc737_f9843783,
        64'hfef42423_2007879b,
        64'h03b907b7_02f71063,
        64'h479d873e_57fcf984,
        64'h3783a275_fef42623,
        64'h47851407_89632781,
        64'hfec42783_fef42623,
        64'h87aa1d40_00eff984,
        64'h35035007_85930319,
        64'h77b7df98_5007071b,
        64'h03197737_f9843783,
        64'hcb2ff0ef_853e0300,
        64'h05934609_43dcf984,
        64'h3783dfc5_27818b89,
        64'hfe442783_aafdfef4,
        64'h26234785_cd6ff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8f984,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_cc4ff0ef,
        64'h853e0300_059343dc,
        64'hf9843783_ac3dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aacbaf_e0eff984,
        64'h35036000_0593863e,
        64'h4681fe84_2783fef4,
        64'h24231007_879b03b9,
        64'h07b70cf7_16634789,
        64'h873e0347_c783f984,
        64'h3783a451_fef42623,
        64'h47852207_85632781,
        64'hfec42783_fef42623,
        64'h87aa2ac0_00eff984,
        64'h350385be_5f9cf984,
        64'h3783df98_0807071b,
        64'h02faf737_f9843783,
        64'hd8aff0ef_853e0300,
        64'h05934609_43dcf984,
        64'h3783dfc5_27818b89,
        64'hfe442783_acd9fef4,
        64'h26234785_daeff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8f984,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_d9cff0ef,
        64'h853e0300_059343dc,
        64'hf9843783_ae19fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aad92f_e0eff984,
        64'h35036000_0593863e,
        64'h4685fe84_2783fef4,
        64'h242337c5_810007b7,
        64'h14e79123_47450000,
        64'h1797fd5f_e0eff984,
        64'h350385be_863afa04,
        64'h07132781_fe245783,
        64'he3aff0ef_853e4591,
        64'h863afe04_570343dc,
        64'hf9843783_fef41023,
        64'h8ff917fd_6785fe04,
        64'h5703fef4_10230400,
        64'h0793fef4_11234785,
        64'hae794785_18e7a923,
        64'h47050000_1797cb3f,
        64'hc0ef2425_05130000,
        64'h151723a5_85930000,
        64'h15971f40_0613a025,
        64'h14f71163_4785873e,
        64'h0347c783_f9843783,
        64'h1c07a223_00001797,
        64'haef94785_1ce7a923,
        64'h47050000_1797cf3f,
        64'hc0ef2825_05130000,
        64'h151727a5_85930000,
        64'h15971f30_0613a025,
        64'h04f71363_11178793,
        64'h111117b7_873e53dc,
        64'hf9843783_2007a423,
        64'h00001797_c385f984,
        64'h3783fc04_3c23fc04,
        64'h3823fc04_3423fc04,
        64'h3023fa04_3c23fa04,
        64'h3823fa04_3423fa04,
        64'h3023f8a4_3c231880,
        64'hf0a2f486_71598082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'he8eff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfc843783_f4eff0ef,
        64'h853e0300_05934609,
        64'h43dcfc84_3783dfc5,
        64'h27818b89_fdc42783,
        64'ha83dfef4_26234785,
        64'hf72ff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fc84_3783c385,
        64'h27818ff9_67a1fdc4,
        64'h2703fcf4_2e2387aa,
        64'hf60ff0ef_853e0300,
        64'h059343dc_fc843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaf56f,
        64'he0effc84_35036000,
        64'h0593863e_4685fe04,
        64'h2783fef4_202337c1,
        64'h010007b7_30e79323,
        64'h47450000_1797998f,
        64'hf0effc84_350385be,
        64'hfc043603_2781fe64,
        64'h5783ffcf_f0ef853e,
        64'h4591863a_fe445703,
        64'h43dcfc84_3783fef4,
        64'h12238ff9_17fd6785,
        64'hfe445703_fef41223,
        64'h04000793_fef41323,
        64'h4785fce7_dee303f0,
        64'h07930007_871bfe84,
        64'h2783fef4_24232785,
        64'hfe842783_00078023,
        64'h97bafc04_3703fe84,
        64'h2783a235_478536e7,
        64'hae234705_00001797,
        64'he9dfc0ef_42c50513,
        64'h00001517_42458593,
        64'h00001597_1a000613,
        64'ha081fe04_24233a07,
        64'ha1230000_1797a285,
        64'h47853ae7_a8234705,
        64'h00001797_ed1fc0ef,
        64'h46050513_00001517,
        64'h45858593_00001597,
        64'h19f00613_a02502f7,
        64'h1d631117_87931111,
        64'h17b7873e_53dcfc84,
        64'h37833e07_a3230000,
        64'h1797c385_fc843783,
        64'hfcb43023_fca43423,
        64'h0080f822_fc067139,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aa851f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783911f,
        64'hf0ef853e_03e00593,
        64'h863a9341_1742fe84,
        64'h270343dc_fd843783,
        64'hfef42423_8fd9fe84,
        64'h278357f8_fd843783,
        64'hfef42423_8ff917e1,
        64'h67c1fe84_2703fef4,
        64'h242387aa_915ff0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_04f71963,
        64'h4791873e_57fcfd84,
        64'h37839edf_f0ef853e,
        64'h02800593_863a0ff7,
        64'h7713fe84_270343dc,
        64'hfd843783_fef42423,
        64'h0027e793_fe842783,
        64'ha039fef4_24230207,
        64'he793fe84_278300f7,
        64'h1963478d_873e0377,
        64'hc783fd84_3783fef4,
        64'h242387aa_9fdff0ef,
        64'h853e0280_059343dc,
        64'hfd843783_8eefd0ef,
        64'h3e800513_9cfff0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe842783,
        64'ha8f5fef4_26234785,
        64'h9f3ff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe84,
        64'h2703fef4_242387aa,
        64'h9e1ff0ef_853e0300,
        64'h059343dc_fd843783,
        64'haa35fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa9d7f,
        64'he0effd84_35036000,
        64'h0593863e_4681fe44,
        64'h2783fef4_22231007,
        64'h879b03b7_07b7a039,
        64'hfef42223_5007879b,
        64'h03b707b7_00f71963,
        64'h4791873e_57fcfd84,
        64'h3783a02d_fef42223,
        64'h2007879b_03b707b7,
        64'ha825fef4_22236007,
        64'h879b03b7_07b700f7,
        64'h19634791_873e57fc,
        64'hfd843783_02f71763,
        64'h478d873e_0377c783,
        64'hfd843783_02e78ba3,
        64'h4709fd84_3783a031,
        64'h02e78ba3_470dfd84,
        64'h378300f7_186347a1,
        64'h873e4bdc_fd843783,
        64'h00f71f63_4795873e,
        64'h0347c783_fd843783,
        64'h02f71763_4789873e,
        64'h0367c783_fd843783,
        64'ha431fef4_26234785,
        64'h12078c63_2781fec4,
        64'h2783fef4_262387aa,
        64'haa9fe0ef_fd843503,
        64'h60078593_67a1863e,
        64'h4681fe44_2783fef4,
        64'h22230377_c783fd84,
        64'h378302e7_8ba34709,
        64'hfd843783_ac81fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaaebf_e0effd84,
        64'h35037007_8593678d,
        64'h863e4681_4bbcfd84,
        64'h378306f7_1b634785,
        64'h873e0347_c783fd84,
        64'h3783a479_fe042623,
        64'h00e7e563_478d873e,
        64'h4bdcfd84_3783a45d,
        64'h47856ae7_ac234705,
        64'h00001797_9d8fd0ef,
        64'h76850513_00001517,
        64'h76058593_00001597,
        64'h11300613_a02504f7,
        64'h10634789_873e0367,
        64'hc783fd84_37836e07,
        64'ha5230000_1797a4dd,
        64'h47856ee7_ac234705,
        64'h00001797_a18fd0ef,
        64'h7a850513_00001517,
        64'h7a058593_00001597,
        64'h11200613_a02504f7,
        64'h13631117_87931111,
        64'h17b7873e_53dcfd84,
        64'h37837207_a7230000,
        64'h1797c385_fd843783,
        64'hfca43c23_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aab95f,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfd84,
        64'h3783c55f_f0ef853e,
        64'h03000593_460943dc,
        64'hfd843783_dfc52781,
        64'h8b89fe04_2783a83d,
        64'hfef42623_4785c79f,
        64'hf0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c3852781,
        64'h8ff967a1_fe042703,
        64'hfef42023_87aac67f,
        64'hf0ef853e_03000593,
        64'h43dcfd84_3783a8bd,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_c5dfe0ef,
        64'hfd843503_30078593,
        64'h67ad4601_86be2781,
        64'hfe645783_80e79323,
        64'h47450000_2797e98f,
        64'hf0effd84_350385be,
        64'hfd043603_2781fe64,
        64'h5783cfdf_f0ef853e,
        64'h4591863a_fe445703,
        64'h43dcfd84_3783fef4,
        64'h12238ff9_17fd6785,
        64'hfe445703_fef41223,
        64'h47a1fef4_13234785,
        64'ha8e5fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aacd7f,
        64'he0effd84_35037007,
        64'h8593678d_863e4681,
        64'h4bbcfd84_3783fce7,
        64'hdfe3479d_0007871b,
        64'hfe842783_fef42423,
        64'h2785fe84_27830007,
        64'h802397ba_fd043703,
        64'hfe842783_aa814785,
        64'h8ae7a323_47050000,
        64'h2797bc6f_d0ef9565,
        64'h05130000_251794e5,
        64'h85930000_25970ba0,
        64'h0613a081_fe042423,
        64'h8c07a623_00002797,
        64'ha2514785_8ce7ad23,
        64'h47050000_2797bfaf,
        64'hd0ef98a5_05130000,
        64'h25179825_85930000,
        64'h25970b90_0613a025,
        64'h02f71d63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_9007a823,
        64'h00002797_c385fd84,
        64'h3783fcb4_3823fca4,
        64'h3c231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_e1fff0ef,
        64'h85364591_863e93c1,
        64'h17c28ff9_17fd6785,
        64'hfd645703_43d4fd84,
        64'h3783fef4_26232781,
        64'h87aad99f_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783a081,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_e05fe0ef,
        64'hfd843503_6585863e,
        64'h46812781_fd645783,
        64'ha0adfef4_26234785,
        64'ha89d4785_9ae7a923,
        64'h47050000_2797cd2f,
        64'hd0efa625_05130000,
        64'h2517a5a5_85930000,
        64'h259707f0_0613a025,
        64'hcb8d2781_3037f793,
        64'hfe842783_fef42423,
        64'h87aae19f_f0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'h9e07ae23_00002797,
        64'ha0f94785_a0e7a523,
        64'h47050000_2797d2af,
        64'hd0efaba5_05130000,
        64'h2517ab25_85930000,
        64'h259707e0_0613a025,
        64'h04f71f63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_a407a023,
        64'h00002797_c385fd84,
        64'h3783fcf4_1b2387ae,
        64'hfca43c23_1800f022,
        64'hf4067179_80826105,
        64'h644260e2_0001eb7f,
        64'hf0ef853e_85bafea4,
        64'h47039381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef40523,
        64'h87bafef4_05a387b6,
        64'hfef42623_873286ae,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e2853e_87aaea9f,
        64'hf0ef853e_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h05a387ba_fef42623,
        64'h872e87aa_1000e822,
        64'hec061101_80826105,
        64'h644260e2_0001f63f,
        64'hf0ef853e_85bafe84,
        64'h57039381_17822781,
        64'h9fb9fec4_27032781,
        64'hfeb44783_fef41423,
        64'h87bafef4_05a387b6,
        64'hfef42623_873286ae,
        64'h87aa1000_e822ec06,
        64'h11018082_61056442,
        64'h60e2853e_87aaf47f,
        64'hf0ef853e_93811782,
        64'h27819fb9_fec42703,
        64'h2781feb4_4783fef4,
        64'h05a387ba_fef42623,
        64'h872e87aa_1000e822,
        64'hec061101_80826145,
        64'h74220001_00e79023,
        64'hfd645703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf41b23_87aefca4,
        64'h3c231800_f4227179,
        64'h80826145_74220001,
        64'h00e78023_fd744703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf40ba3,
        64'h87aefca4_3c231800,
        64'hf4227179_80826105,
        64'h6462853e_2781439c,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61056462_853e93c1,
        64'h17c20007_d783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826105,
        64'h6462853e_0ff7f793,
        64'h0007c783_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61616406,
        64'h60a6853e_fec42783,
        64'hfe042623_d3f8fb84,
        64'h37830007_871b0097,
        64'hd79bfd84_2783fcf4,
        64'h2c2302f7_07bbfe04,
        64'h2783fd84_2703fcf4,
        64'h2c2302f7_07bbfdc4,
        64'h27032781_2785fd84,
        64'h2783fcf4_2c238fd9,
        64'hfd842783_0007871b,
        64'h8ff9c007_87936785,
        64'h873e2781_00a7979b,
        64'hfd042783_fcf42c23,
        64'h0167d79b_fcc42783,
        64'hfcf42e23_278100f7,
        64'h17bb4705_27812789,
        64'h27818b9d_27810077,
        64'hd79bfcc4_2783fef4,
        64'h20232781_00f717bb,
        64'h47052781_8bbd2781,
        64'h0087d79b_fd042783,
        64'h02e78aa3_fb843783,
        64'h0ff7f713_8bbd0ff7,
        64'hf7932781_0127d79b,
        64'hfd442783_fcf42a23,
        64'h278187aa_9bdfd0ef,
        64'h853e9381_17822781,
        64'h27f143dc_fb843783,
        64'hfcf42823_278187aa,
        64'h9d9fd0ef_853e9381,
        64'h17822781_27e143dc,
        64'hfb843783_fcf42623,
        64'h278187aa_9f5fd0ef,
        64'h853e9381_17822781,
        64'h27d143dc_fb843783,
        64'hfcf42423_278187aa,
        64'ha11fd0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_a23dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa9d2f_f0effb84,
        64'h35039007_85936785,
        64'h863e4681_4bbcfb84,
        64'h3783aab1_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'ha00ff0ef_fb843503,
        64'h30000593_863e4681,
        64'h4bbcfb84_3783cbb8,
        64'h12340737_fb843783,
        64'hc7f8fb84_37830007,
        64'h871b87aa_b31fd0ef,
        64'h853e45f1_43dcfb84,
        64'h3783c7b8_fb843783,
        64'h0007871b_87aab4bf,
        64'hd0ef853e_45e143dc,
        64'hfb843783_c3f8fb84,
        64'h37830007_871b87aa,
        64'hb65fd0ef_853e45d1,
        64'h43dcfb84_3783c3b8,
        64'hfb843783_0007871b,
        64'h87aab7ff_d0ef853e,
        64'h45c143dc_fb843783,
        64'haaedfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaa9ef,
        64'hf0effb84_35032000,
        64'h05934601_4681db98,
        64'h4705fb84_3783c789,
        64'h27818ff9_400007b7,
        64'hfe842703_fa07dde3,
        64'hfe842783_fef42423,
        64'h87aab3bf_d0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783aca1,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_afcff0ef,
        64'hfb843503_10000593,
        64'h40ff8637_4681a091,
        64'hfe042423_a459fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aab2af_f0effb84,
        64'h35034581_46014681,
        64'ha46dfef4_26234785,
        64'he7892781_8ff967c1,
        64'hfe442703_fef42223,
        64'h87aabbbf_d0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fb843783,
        64'hcb8d47dc_fb843783,
        64'h02f70e63_400007b7,
        64'h873e2781_8ff9c000,
        64'h07b7873e_579cfb84,
        64'h3783a601_4785f0e7,
        64'hae234705_00002797,
        64'ha3dfd0ef_fac50513,
        64'h00002517_fac58593,
        64'h00002597_67100613,
        64'ha02504f7_13634789,
        64'h873e0367_c783fb84,
        64'h3783f407_a7230000,
        64'h2797a681_4785f4e7,
        64'hae234705_00002797,
        64'ha7dfd0ef_fec50513,
        64'h00002517_fec58593,
        64'h00002597_67000613,
        64'ha02504f7_13631117,
        64'h87931111_17b7873e,
        64'h53dcfb84_3783f807,
        64'ha9230000_2797c385,
        64'hfb843783_faa43c23,
        64'h0880e0a2_e486715d,
        64'h80826121_744270e2,
        64'h0001d05f_d0ef853a,
        64'h85be2781_08078793,
        64'hfd843783_93010207,
        64'h97132781_0587879b,
        64'h43dcfd84_378300e7,
        64'h912397b6_078e07c1,
        64'h93810206_1793fd84,
        64'h36839341_03079713,
        64'h02f707bb_0006861b,
        64'h36fdfec4_268393c1,
        64'h17c2fe44_27839341,
        64'h03079713_fd442783,
        64'h00e79023_02300713,
        64'h97ba078e_07c19381,
        64'h1782fd84_37032781,
        64'h37fdfec4_2783c3d8,
        64'h97b6078e_07c19381,
        64'h02061793_fd843683,
        64'h0007871b_9fb90006,
        64'h861b36fd_fec42683,
        64'h27810107_979bfe84,
        64'h27830007_871bfc84,
        64'h3783f8e7_ebe32781,
        64'hfe842783_0007871b,
        64'h37fdfec4_2783fef4,
        64'h24232785_fe842783,
        64'h00079123_97ba078e,
        64'h07c1fe84_6783fd84,
        64'h370300e7_90230210,
        64'h071397ba_078e07c1,
        64'hfe846783_fd843703,
        64'hc3d897b6_078e07c1,
        64'hfe846783_fd843683,
        64'h0007871b_9fb92781,
        64'h0107979b_fe842783,
        64'h0007871b_fc843783,
        64'ha8b1fe04_2423fef4,
        64'h26232785_fec42783,
        64'hc7912781_8ff917fd,
        64'h67c1873e_278102f7,
        64'h07bbfe44_2783fd44,
        64'h2703fef4_26230107,
        64'hd79b2781_02f707bb,
        64'hfe442783_fd442703,
        64'ha835fef4_26234785,
        64'h00f77663_67c1873e,
        64'h278102f7_07bbfe44,
        64'h2783fd44_2703fef4,
        64'h22238ff9_17fd6785,
        64'hfe442703_fef42223,
        64'h87aaebff_d0ef853e,
        64'h459143dc_fd843783,
        64'hfe042223_fe042423,
        64'hfe042623_fcf42a23,
        64'hfcc43423_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_61457402,
        64'h70a2853e_fec42783,
        64'h0001a011_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'he10ff0ef_fd843503,
        64'h70000593_863e4681,
        64'h4bbcfd84_3783fe04,
        64'h2623fca4_3c231800,
        64'hf022f406_71798082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hf87fd0ef_853e0300,
        64'h05934609_43dcfd84,
        64'h3783dfc5_27818b89,
        64'hfe442783_a00dfef4,
        64'h26234785_fabfd0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_f99fd0ef,
        64'h853e0300_059343dc,
        64'hfd843783_a08dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaebaf_f0effd84,
        64'h35039007_85936789,
        64'h863e86ba_fd442783,
        64'hfd042703_26e79423,
        64'h02700713_00002797,
        64'ha879fef4_26234785,
        64'hc3b92781_fec42783,
        64'hfef42623_87aaef6f,
        64'hf0effd84_35038007,
        64'h85936789_863e86ba,
        64'hfd442783_fd042703,
        64'h2ae79123_470d0000,
        64'h279702f7_1f634785,
        64'h0007871b_fd042783,
        64'h142000ef_fd843503,
        64'h85befc84_3603fd04,
        64'h2783a8e5_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h081000ef_fd843503,
        64'h20000593_02f70363,
        64'h20000793_873e2781,
        64'h87aafd3f_d0ef853e,
        64'h93811782_27812791,
        64'h43dcfd84_3783aa35,
        64'hfef42623_4785e789,
        64'h27818ff9_67c1fe84,
        64'h2703fef4_242387aa,
        64'h800fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783cb8d,
        64'h47dcfd84_378302f7,
        64'h0e634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_fd843783,
        64'h00f71f63_4789873e,
        64'h0367c783_fd843783,
        64'hfcf42823_87bafcf4,
        64'h2a23fcd4_34238732,
        64'h87aefca4_3c230080,
        64'hf822fc06_71398082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'h880fe0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfd843783_96afe0ef,
        64'h853e0300_05934609,
        64'h43dcfd84_3783dfc5,
        64'h27818b89_fe442783,
        64'ha83dfef4_26234785,
        64'h98efe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783c385,
        64'h27818ff9_67a1fe44,
        64'h2703fef4_222387aa,
        64'h97cfe0ef_853e0300,
        64'h059343dc_fd843783,
        64'ha8bdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa89ff,
        64'hf0effd84_35032007,
        64'h85936785_863e86ba,
        64'hfd442783_fd042703,
        64'h44e79623_03700713,
        64'h00002797_a86dfef4,
        64'h26234785_c3b92781,
        64'hfec42783_fef42623,
        64'h87aa8dbf_f0effd84,
        64'h35031007_85936785,
        64'h863e86ba_fd442783,
        64'hfd042703_48e79323,
        64'h474d0000_279702f7,
        64'h1f634785_0007871b,
        64'hfd042783_326000ef,
        64'hfd843503_85befc84,
        64'h3603fd04_2783aa11,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_265000ef,
        64'hfd843503_20000593,
        64'h02f70363_20000793,
        64'h873e2781_87aa9b6f,
        64'he0ef853e_93811782,
        64'h27812791_43dcfd84,
        64'h3783aaa1_fef42623,
        64'h4785e789_27818ff9,
        64'h67c1fe84_2703fef4,
        64'h242387aa_9e4fe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783cb8d_47dcfd84,
        64'h378302f7_0e634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfd843783_00f71f63,
        64'h4789873e_0367c783,
        64'hfd843783_fcf42823,
        64'h87bafcf4_2a23fcd4,
        64'h34238732_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_61457422,
        64'h853efec4_27830001,
        64'ha0110001_a0210001,
        64'ha031fef4_26238fd9,
        64'hfd442783_fec42703,
        64'ha831fef4_262301a7,
        64'he793fec4_2783a02d,
        64'hfef42623_03a7e793,
        64'hfec42783_a825fef4,
        64'h262301a7_e793fec4,
        64'h2783a099_fef42623,
        64'h0027e793_fec42783,
        64'ha891fef4_262303a7,
        64'he793fec4_2783a08d,
        64'hfef42623_03a7e793,
        64'hfec42783_a885fef4,
        64'h262301a7_e793fec4,
        64'h2783a8bd_fef42623,
        64'h0097e793_fec42783,
        64'ha071fef4_262303a7,
        64'he793fec4_2783a869,
        64'hfef42623_01a7e793,
        64'hfec42783_00f71963,
        64'h4785873e_0347c783,
        64'hfd843783_a865fef4,
        64'h262301a7_e793fec4,
        64'h2783a0d9_fef42623,
        64'h01a7e793_fec42783,
        64'ha8d1fef4_262301b7,
        64'he793fec4_2783a0cd,
        64'hfef42623_03a7e793,
        64'hfec42783_00f71963,
        64'h4785873e_0347c783,
        64'hfd843783_a201fef4,
        64'h262301b7_e793fec4,
        64'h2783a239_fef42623,
        64'h01b7e793_fec42783,
        64'haa31fef4_26230097,
        64'he793fec4_2783a22d,
        64'hfef42623_0027e793,
        64'hfec42783_aa390ef7,
        64'h05639007_879367ad,
        64'h0007871b_10e68a63,
        64'h30070713_672d0007,
        64'h869b10e6_8a63a007,
        64'h0713672d_0007869b,
        64'ha2a916f7_0363a007,
        64'h87936791_0007871b,
        64'h0ee68d63_d0070713,
        64'h67250007_869b0ae6,
        64'h89636007_07136721,
        64'h0007869b_02d76863,
        64'h70070713_67250007,
        64'h869b14e6_80637007,
        64'h07136725_0007869b,
        64'haa4914f7_08638007,
        64'h87936789_0007871b,
        64'h18e68b63_40070713,
        64'h670d0007_869b16e6,
        64'h86639007_07136709,
        64'h0007869b_aa7d16f7,
        64'h07632007_87936785,
        64'h0007871b_16e68e63,
        64'h50070713_67050007,
        64'h869b18e6_85633007,
        64'h07136705_0007869b,
        64'h02d76863_70070713,
        64'h67050007_869b1ae6,
        64'h8a637007_07136705,
        64'h0007869b_06d76c63,
        64'h70070713_670d0007,
        64'h869b20e6_84637007,
        64'h0713670d_0007869b,
        64'ha40d1cf7_0263b007,
        64'h87936785_0007871b,
        64'h1ce68963_67050007,
        64'h869b1ce6_8e63c007,
        64'h07136705_0007869b,
        64'ha4a91af7_02637000,
        64'h07930007_871b1ee6,
        64'h85639007_07136705,
        64'h0007869b_1c070663,
        64'h27018007_871b02d7,
        64'h6563a007_07136705,
        64'h0007869b_20e68f63,
        64'ha0070713_67050007,
        64'h869ba471_18f70863,
        64'h30000793_0007871b,
        64'h1ae68563_50000713,
        64'h0007869b_2ae68e63,
        64'h40000713_0007869b,
        64'hac4d18f7_0d631000,
        64'h07930007_871b2c07,
        64'h09630007_871b00d7,
        64'h6d632000_07130007,
        64'h869b1ce6_84632000,
        64'h07130007_869b04d7,
        64'h6c636000_07130007,
        64'h869b20e6_85636000,
        64'h07130007_869b0cd7,
        64'h6d631007_07136705,
        64'h0007869b_2ae68a63,
        64'h10070713_67050007,
        64'h869bfd44_2783fef4,
        64'h2623fd44_2783fcf4,
        64'h2a2387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'he86fe0ef_853e0300,
        64'h05934605_43dcfd84,
        64'h3783d3a9_27818b85,
        64'hfe042783_a00dea4f,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_fef42623,
        64'h4789e781_27819bf9,
        64'hfec42783_fef42623,
        64'h87aae96f_e0ef853e,
        64'h03200593_43dcfd84,
        64'h3783c3a1_27818ff9,
        64'h67a1fe04_2703a899,
        64'heeefe0ef_853e0300,
        64'h05930200_061343dc,
        64'hfd843783_cf812781,
        64'h0207f793_278187aa,
        64'hed4fe0ef_853e0300,
        64'h059343dc_fd843783,
        64'h02f71b63_30078793,
        64'h67850007_871bfd44,
        64'h278300f7_0b635007,
        64'h87936785_0007871b,
        64'hfd442783_fef42023,
        64'h87aaf0ef_e0ef853e,
        64'h03000593_43dcfd84,
        64'h3783ef4f_e0ef853a,
        64'h85be2781_8fd52781,
        64'h9b87d783_00003797,
        64'h0007869b_0107979b,
        64'hfe442783_93010207,
        64'h97132781_27b143dc,
        64'hfd843783_a229fef4,
        64'h26234785_c7892781,
        64'h0207f793_fe442783,
        64'hcb992781_8b89fe84,
        64'h2783fef4_242387aa,
        64'hed8fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_378302f7,
        64'h0f633007_87936785,
        64'h0007871b_fd442783,
        64'h04f70863_50078793,
        64'h67850007_871bfd44,
        64'h2783fef4_22238ff9,
        64'h17fd6791_fe442703,
        64'hfef42223_87aa18c0,
        64'h00effd84_350385be,
        64'hfd442783_80bfe0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783821f_e0ef853a,
        64'h03000593_fff78613,
        64'h67c143d8_fd843783,
        64'hfd2fe0ef_853e85ba,
        64'hfd042703_93811782,
        64'h278127a1_43dcfd84,
        64'h37838d1f_e0ef853e,
        64'h02e00593_463943dc,
        64'hfd843783_863fe0ef,
        64'h853e4599_863a9341,
        64'h1742fcc4_270343dc,
        64'hfd843783_aaedfef4,
        64'h26234785_a4194785,
        64'hace7ab23_47050000,
        64'h3797df6f_e0efb665,
        64'h05130000_3517b665,
        64'h85930000_359744c0,
        64'h0613a025_cb8d2781,
        64'h8b85fe84_2783fef4,
        64'h242387aa_fe4fe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783b007_af230000,
        64'h3797acb1_4785b2e7,
        64'ha6234705_00003797,
        64'he4cfe0ef_bbc50513,
        64'h00003517_bbc58593,
        64'h00003597_44b00613,
        64'ha02504f7_1e631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783b607,
        64'ha1230000_3797c385,
        64'hfd843783_fcf42623,
        64'h87bafcf4_282387b2,
        64'hfcf42a23_873687ae,
        64'hfca43c23_0080f822,
        64'hfc067139_80826145,
        64'h740270a2_853efec4,
        64'h27830001_fcf719e3,
        64'h01f007b7_873e2781,
        64'h8ff901f0_07b7fe84,
        64'h2703fef4_242387aa,
        64'h899fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783a839,
        64'hfef42423_87aa8b7f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_ff6fe0ef,
        64'h3e800513_9abfe0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0047e793,
        64'h93c117c2_fe442783,
        64'h43d8fd84_3783fef4,
        64'h222387aa_999fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_d3ed2781,
        64'h8b89fe44_2783fef4,
        64'h222387aa_9b9fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a821fef4,
        64'h222387aa_9d1fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a1bfe0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0017e793,
        64'h93c117c2_fe442783,
        64'h43d8fd84_3783fef4,
        64'h222387aa_a09fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a211fef4,
        64'h26234785_e7892781,
        64'h8ba12781_fe245783,
        64'hfef41123_87aaa33f,
        64'he0ef853e_03e00593,
        64'h43dcfd84_37838d1f,
        64'he0ef3887_85136785,
        64'ha87fe0ef_853e03e0,
        64'h0593863a_fe245703,
        64'h43dcfd84_3783fef4,
        64'h11230087_e793fe24,
        64'h5783fef4_112387aa,
        64'ha75fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'habffe0ef_853e02c0,
        64'h0593863a_fe245703,
        64'h43dcfd84_3783fef4,
        64'h11239be9_fe245783,
        64'hfef41123_87aaaabf,
        64'he0ef853e_02c00593,
        64'h43dcfd84_3783ffe1,
        64'h27818ff9_01f007b7,
        64'hfe842703_fef42423,
        64'h87aaa33f_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'ha839fef4_242387aa,
        64'ha51fe0ef_853e9381,
        64'h17822781_0247879b,
        64'h43dcfd84_3783fef4,
        64'h26234785_c7812781,
        64'hfec42783_fef42623,
        64'h87aa2120_00effd84,
        64'h3503b007_85936785,
        64'h46014681_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623f3e5_27818b89,
        64'h2781feb4_4783fef4,
        64'h05a387aa_bd9fe0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_a821fef4,
        64'h05a387aa_bf1fe0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_c3bfe0ef,
        64'h853e02f0_05934609,
        64'h43dcfd84_3783bcdf,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_be3fe0ef,
        64'h853a0300_0593fff7,
        64'h861367c1_43d8fd84,
        64'h378302e7_8a234709,
        64'hfd843783_a03102e7,
        64'h8a234705_fd843783,
        64'hc7992781_fec42783,
        64'hfef42623_87aa2de0,
        64'h00effd84_35031000,
        64'h059340ff_86374681,
        64'ha855fef4_26234785,
        64'ha0c14785_e8e7a523,
        64'h47050000_37979abf,
        64'he0eff1a5_05130000,
        64'h3517f1a5_85930000,
        64'h35973ac0_0613a025,
        64'hcb8d2781_fec42783,
        64'hfef42623_87aa32e0,
        64'h00effd84_35034581,
        64'h46014681_acffe0ef,
        64'h71078513_6789ec07,
        64'ha9230000_3797aa19,
        64'h4785eee7_a0234705,
        64'h00003797_a01fe0ef,
        64'hf7050513_00003517,
        64'hf7058593_00003597,
        64'h3ab00613_a02504f7,
        64'h1e631117_87931111,
        64'h17b7873e_53dcfd84,
        64'h3783f007_ab230000,
        64'h3797c385_fd843783,
        64'hfca43c23_1800f022,
        64'hf4067179_8082614d,
        64'h64ea740a_70aa853e,
        64'hfdc42783_0001a011,
        64'h0001a021_0001a031,
        64'hfcf42e23_4785cb89,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_504010ef,
        64'hf5843503_20000593,
        64'h02f71763_4785873e,
        64'h0347c783_f5843783,
        64'h00f71a63_4791873e,
        64'h57fcf584_37830001,
        64'ha0b9fcf4_2e234785,
        64'hc7912781_fdc42783,
        64'hfcf42e23_87aa79e0,
        64'h20eff584_350385be,
        64'hfd442783_fcf42a23,
        64'h1007879b_03a207b7,
        64'heb950a27_c783dbe7,
        64'h87930000_3797a071,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_09d010ef,
        64'hf5843503_02f71163,
        64'h4791873e_57fcf584,
        64'h3783a865_fcf42e23,
        64'h478500f7_06634785,
        64'h873e0b97_c783e067,
        64'h87930000_379704f7,
        64'h16634791_873e57fc,
        64'hf5843783_00f70963,
        64'h4795873e_57fcf584,
        64'h3783a8c5_fcf42e23,
        64'h478500f7_06634789,
        64'h873e0b97_c783e3e7,
        64'h87930000_379702f7,
        64'h1063479d_873e57fc,
        64'hf5843783_aa29fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa6ac0_20eff584,
        64'h3503e725_85930000,
        64'h3597a281_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h657010ef_f5843503,
        64'h0cf70b63_4799873e,
        64'h57fcf584_3783d7f8,
        64'h4719f584_3783a029,
        64'hd7f84715_f5843783,
        64'h00e7f763_4785873e,
        64'h0377c783_f5843783,
        64'hcf912781_8b892781,
        64'h0c47c783_ed478793,
        64'h00003797_a825d7f8,
        64'h4711f584_378300e7,
        64'hf7634785_873e0377,
        64'hc783f584_3783cf91,
        64'h27818bb1_27810c47,
        64'hc783f027_87930000,
        64'h3797a09d_d7f8471d,
        64'hf5843783_00e7f763,
        64'h4785873e_0377c783,
        64'hf5843783_cf912781,
        64'h0307f793_27810c47,
        64'hc783f327_87930000,
        64'h3797d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0d47c783_f4c78793,
        64'h00003797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0087979b_27810d57,
        64'hc783f727_87930000,
        64'h379753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810107,
        64'h979b2781_0d67c783,
        64'hf9878793_00003797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h0187979b_27810d77,
        64'hc783fba7_87930000,
        64'h3797a461_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h01b020ef_f5843503,
        64'hfe058593_00003597,
        64'ha47dfcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa2bf0,
        64'h10eff584_350328f7,
        64'h12634795_873e0347,
        64'hc783f584_3783acf1,
        64'hfcf42e23_478528f7,
        64'h0d634785_873e0b97,
        64'hc78302a7_87930000,
        64'h3797ace5_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h08b020ef_f5843503,
        64'h05058593_00003597,
        64'hae39fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa0340,
        64'h20eff584_3503d7f8,
        64'h4715f584_37832ee7,
        64'hfd634785_873e0377,
        64'hc783f584_37833007,
        64'h85632781_8b892781,
        64'h0c47c783_09c78793,
        64'h00003797_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810d47_c7830b67,
        64'h87930000_379753f8,
        64'hf5843783_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810087_979b2781,
        64'h0d57c783_0dc78793,
        64'h00003797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_8fd92781,
        64'h0107979b_27810d67,
        64'hc7831027_87930000,
        64'h379753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b0187_979b2781,
        64'h0d77c783_12478793,
        64'h00003797_aecdfcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa1850_20eff584,
        64'h350314a5_85930000,
        64'h3597a921_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h429010ef_f5843503,
        64'h14f71f63_4785873e,
        64'h0367c783_f5843783,
        64'h16e7f763_478d873e,
        64'h0357c783_f5843783,
        64'h16f71f63_4789873e,
        64'h0347c783_f5843783,
        64'ha19dfcf4_2e234785,
        64'h42078363_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h17e020ef_f5843503,
        64'hd7f84715_f5843783,
        64'h44e7f363_4785873e,
        64'h0377c783_f5843783,
        64'h44078b63_27818b89,
        64'h2781f9d4_47834607,
        64'h82630004_c78302e7,
        64'h8e234705_f5843783,
        64'h802ff0ef_3e800513,
        64'h9b6ff0ef_853a02c0,
        64'h0593863e_93c117c2,
        64'h0047e793_fda45783,
        64'h43d8f584_3783fcf4,
        64'h1d2387aa_9a0ff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_d3e52781,
        64'h8b892781_fda45783,
        64'hfcf41d23_87aa9c2f,
        64'hf0ef853e_02c00593,
        64'h43dcf584_3783a821,
        64'hfcf41d23_87aa9daf,
        64'hf0ef853e_02c00593,
        64'h43dcf584_3783a24f,
        64'hf0ef853a_02c00593,
        64'h863e93c1_17c20017,
        64'he793fda4_578343d8,
        64'hf5843783_fcf41d23,
        64'h87aaa0ef_f0ef853e,
        64'h02c00593_43dcf584,
        64'h3783a3a5_fcf42e23,
        64'h4785e789_27818ba1,
        64'h2781fd24_5783fcf4,
        64'h192387aa_a38ff0ef,
        64'h853e03e0_059343dc,
        64'hf5843783_8d6ff0ef,
        64'h38878513_6785a8cf,
        64'hf0ef853e_03e00593,
        64'h863afd24_570343dc,
        64'hf5843783_fcf41923,
        64'h0087e793_fd245783,
        64'hfcf41923_87aaa7af,
        64'hf0ef853e_03e00593,
        64'h43dcf584_3783ac4f,
        64'hf0ef853e_02c00593,
        64'h863afd24_570343dc,
        64'hf5843783_fcf41923,
        64'h9be9fd24_5783fcf4,
        64'h192387aa_ab0ff0ef,
        64'h853e02c0_059343dc,
        64'hf5843783_14079d63,
        64'h03c7c783_f5843783,
        64'h16f71363_47a1873e,
        64'h4bdcf584_378316e7,
        64'hfa63478d_873ef9d4,
        64'h47831807_d0634187,
        64'hd79b0187_979b0024,
        64'hc7836207_9e632781,
        64'hfdc42783_fcf42e23,
        64'h87aa18e0_20eff584,
        64'h350385be_f9040793,
        64'hadb9fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa66f0,
        64'h10eff584_3503c385,
        64'h27818b91_27810014,
        64'hc783a561_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h4b3010ef_f5843503,
        64'h85a6a565_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h34d020ef_f5843503,
        64'h26f71263_4785873e,
        64'h0347c783_f5843783,
        64'hadd9fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa46c0,
        64'h10eff584_3503add5,
        64'hfcf42e23_4785adf5,
        64'hfcf42e23_4785cb89,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_06f020ef,
        64'hf5843503_85be5f9c,
        64'hf5843783_df98a807,
        64'h071b018c_c737f584,
        64'h3783af05_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h6dc010ef_f5843503,
        64'h04f71b63_4795873e,
        64'h0347c783_f5843783,
        64'h00f70a63_4789873e,
        64'h0347c783_f5843783,
        64'ha7bdfcf4_2e234785,
        64'hc3d12781_fdc42783,
        64'hfcf42e23_87aa0e10,
        64'h20eff584_350385be,
        64'h5f9cf584_3783df98,
        64'h8407071b_017d8737,
        64'hf5843783_a801df98,
        64'hac07071b_0121f737,
        64'hf5843783_00f71a63,
        64'h4789873e_0367c783,
        64'hf5843783_7c40006f,
        64'hfcf42e23_4785c791,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_915ff0ef,
        64'hf5843503_06f71c63,
        64'h4785873e_0347c783,
        64'hf5843783_7f40006f,
        64'hfcf42e23_478500f7,
        64'h07634795_873e0347,
        64'hc783f584_378300f7,
        64'h0f634789_873e0347,
        64'hc783f584_378302f7,
        64'h07634785_873e0347,
        64'hc783f584_378302f7,
        64'h02e34785_0007871b,
        64'hfdc42783_fcf42e23,
        64'h87aa0530_00eff584,
        64'h3503a839_02e78a23,
        64'h4715f584_378300f7,
        64'h18634000_07b7873e,
        64'h27818ff9_c00007b7,
        64'h873e579c_f5843783,
        64'h0750006f_47857ae7,
        64'haa234705_00003797,
        64'had4ff0ef_84450513,
        64'h00004517_84458593,
        64'h00004597_24000613,
        64'ha02d04f7_1a634789,
        64'h873e0367_c783f584,
        64'h3783df98_a807071b,
        64'h00062737_f5843783,
        64'h02078e23_f5843783,
        64'h02e78a23_4705f584,
        64'h378302e7_8ba34705,
        64'hf5843783_8007a823,
        64'h00004797_0e10006f,
        64'h478582e7_a0234705,
        64'h00004797_b40ff0ef,
        64'h8b050513_00004517,
        64'h8b058593_00004597,
        64'h23f00613_a02d06f7,
        64'h19631117_87931111,
        64'h17b7873e_53dcf584,
        64'h37838407_ab230000,
        64'h4797c385_f5843783,
        64'hfc043423_fc043023,
        64'hfa043c23_fa043823,
        64'hfa043423_fa043023,
        64'hf8043c23_f8043823,
        64'h0004b023_00579493,
        64'h839507fd_f8078793,
        64'hfe040793_f4a43c23,
        64'h1900ed26_f122f506,
        64'h71718082_61616406,
        64'h60a6853e_fec42783,
        64'hfe042623_d3f8fb84,
        64'h37830007_871b00a7,
        64'h979b2781_27852781,
        64'h8ff917fd_004007b7,
        64'h873e2781_0087d79b,
        64'hfc442783_02f71663,
        64'h4785873e_27818b8d,
        64'h27810167_d79bfcc4,
        64'h2783a081_d3f8fb84,
        64'h37830007_871b0097,
        64'hd79bfd04_2783fcf4,
        64'h282302f7_07bbfd84,
        64'h2783fd04_2703fcf4,
        64'h282302f7_07bbfd44,
        64'h27032781_2785fd04,
        64'h2783fcf4_28238fd9,
        64'hfd042783_0007871b,
        64'h8ff9c007_87936785,
        64'h873e2781_00a7979b,
        64'hfc842783_fcf42823,
        64'h0167d79b_fc442783,
        64'hfcf42a23_278100f7,
        64'h17bb4705_27812789,
        64'h27818b9d_27810077,
        64'hd79bfc44_2783fcf4,
        64'h2c232781_00f717bb,
        64'h47052781_8bbd2781,
        64'h0087d79b_fc842783,
        64'he3c52781_8b8d2781,
        64'h0167d79b_fcc42783,
        64'hfcf42623_278187aa,
        64'he88ff0ef_853e9381,
        64'h17822781_27f143dc,
        64'hfb843783_fcf42423,
        64'h278187aa_ea4ff0ef,
        64'h853e9381_17822781,
        64'h27e143dc_fb843783,
        64'hfcf42223_278187aa,
        64'hec0ff0ef_853e9381,
        64'h17822781_27d143dc,
        64'hfb843783_fcf42023,
        64'h278187aa_edcff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'ha28dfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa69f0,
        64'h00effb84_35039007,
        64'h85936785_863e4681,
        64'h4bbcfb84_3783d7d5,
        64'h4bbcfb84_3783cbb8,
        64'hfb843783_0007871b,
        64'h8ff977c1_873e2781,
        64'h87aaf3af_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783a2c1,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_6fd000ef,
        64'hfb843503_30000593,
        64'h46014681_c7f8fb84,
        64'h37830007_871b87aa,
        64'h81dff0ef_853e45f1,
        64'h43dcfb84_3783c7b8,
        64'hfb843783_0007871b,
        64'h87aa837f_f0ef853e,
        64'h45e143dc_fb843783,
        64'hc3f8fb84_37830007,
        64'h871b87aa_851ff0ef,
        64'h853e45d1_43dcfb84,
        64'h3783c3b8_fb843783,
        64'h0007871b_87aa86bf,
        64'hf0ef853e_45c143dc,
        64'hfb843783_a4b9fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa78b0_00effb84,
        64'h35032000_05934601,
        64'h4681ac95_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h585000ef_fb843503,
        64'h02e78e23_4705fb84,
        64'h3783c78d_27818ff9,
        64'h010007b7_fe842703,
        64'hdb984705_fb843783,
        64'hc7892781_8ff94000,
        64'h07b7fe84_2703f407,
        64'hdde3fe84_2783fef4,
        64'h242387aa_85dff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'ha4cdfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa01e0,
        64'h10effb84_35039007,
        64'h859367ad_863e4681,
        64'hfe442783_fef42223,
        64'h8fd90100_07b7fe44,
        64'h270300f7_196347a1,
        64'h873e4bdc_fb843783,
        64'h02f71063_4789873e,
        64'h0367c783_fb843783,
        64'hfef42223_40ff87b7,
        64'ha689fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa07e0,
        64'h10effb84_35037007,
        64'h8593678d_46014681,
        64'ha055fe04_242302e7,
        64'h8aa34709_fb843783,
        64'ha03102e7_8aa34705,
        64'hfb843783_00f70863,
        64'h1aa00793_0007871b,
        64'hfe842783_fef42423,
        64'h87aa92bf_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfb84_3783f3e5,
        64'h27818b89_2781fe34,
        64'h4783fef4_01a387aa,
        64'ha6dff0ef_853e02f0,
        64'h059343dc_fb843783,
        64'ha821fef4_01a387aa,
        64'ha85ff0ef_853e02f0,
        64'h059343dc_fb843783,
        64'hacfff0ef_853e02f0,
        64'h05934609_43dcfb84,
        64'h378304f7_18634789,
        64'h0007871b_fec42783,
        64'ha129fef4_26234785,
        64'h00f70663_47890007,
        64'h871bfec4_2783cf81,
        64'h2781fec4_2783fef4,
        64'h262387aa_154010ef,
        64'hfb843503_80078593,
        64'h67851aa0_06134681,
        64'ha189fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa17e0,
        64'h10effb84_35034581,
        64'h46014681_a19dfef4,
        64'h26234785_e7892781,
        64'h8ff967c1_fdc42703,
        64'hfcf42e23_87aaa0ff,
        64'hf0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfb843783_cb8d47dc,
        64'hfb843783_02f70e63,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cfb84_3783a975,
        64'h4785d6e7_a8234705,
        64'h00004797_891ff0ef,
        64'he0050513_00004517,
        64'he0058593_00004597,
        64'h16200613_a02504f7,
        64'h13634789_873e0367,
        64'hc783fb84_3783cbd8,
        64'h4711fb84_3783da07,
        64'ha5230000_4797a311,
        64'h4785dae7_ac234705,
        64'h00004797_8d9ff0ef,
        64'he4850513_00004517,
        64'he4858593_00004597,
        64'h16100613_a02504f7,
        64'h17631117_87931111,
        64'h17b7873e_53dcfb84,
        64'h3783de07_a7230000,
        64'h4797c385_fb843783,
        64'hfaa43c23_0880e0a2,
        64'he486715d_80826121,
        64'h744270e2_853efec4,
        64'h2783fe04_2623bcdf,
        64'hf0ef853e_45912000,
        64'h061343dc_fd843783,
        64'he2e79923_474d0000,
        64'h4797be9f_f0ef853e,
        64'h03a00593_460143dc,
        64'hfd843783_bfbff0ef,
        64'h853e0380_05934601,
        64'h43dcfd84_3783c0df,
        64'hf0ef853a_03600593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c23ff0ef,
        64'h853a0340_0593eff7,
        64'h861367c1_43d8fd84,
        64'h3783cb9f_f0ef853e,
        64'h02800593_464143dc,
        64'hfd843783_ccbff0ef,
        64'h853a0290_0593863e,
        64'h0ff7f793_0017e793,
        64'hfeb44783_43d8fd84,
        64'h3783fe04_05a3a019,
        64'hfef405a3_47a9c789,
        64'h27818ff9_040007b7,
        64'h873e579c_fd843783,
        64'ha005fef4_05a347b1,
        64'hc7892781_8ff90200,
        64'h07b7873e_579cfd84,
        64'h3783a82d_fef405a3,
        64'h47b9c789_27818ff9,
        64'h010007b7_873e579c,
        64'hfd843783_a8d5fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa13c0_30effd84,
        64'h3503a807_85930006,
        64'h27b7b35f_f0ef0c80,
        64'h051300f7_16634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfd843783_02f71363,
        64'h4789873e_0367c783,
        64'hfd843783_d93ff0ef,
        64'h853e0290_0593463d,
        64'h43dcfd84_3783a811,
        64'hda7ff0ef_853e0290,
        64'h0593463d_43dcfd84,
        64'h378300f7_1c634789,
        64'h873e0367_c783fd84,
        64'h3783d798_fd843783,
        64'h0007871b_87aac7ff,
        64'hf0ef853e_93811782,
        64'h27810407_879b43dc,
        64'hfd843783_02e78b23,
        64'hfd843783_0ff7f713,
        64'h87aad3ff_f0ef853e,
        64'h0fe00593_43dcfd84,
        64'h3783f3e5_27818b85,
        64'h2781fea4_4783fef4,
        64'h052387aa_de1ff0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_a821fef4,
        64'h052387aa_df9ff0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_e43ff0ef,
        64'h853e02f0_05934605,
        64'h43dcfd84_3783c29f,
        64'hf0ef3e80_0513e5df,
        64'hf0ef853e_02900593,
        64'h460143dc_fd843783,
        64'ha811e71f_f0ef853e,
        64'h02900593_464143dc,
        64'hfd843783_a4814785,
        64'h04e7ab23_47050000,
        64'h4797b77f_f0ef0e65,
        64'h05130000_45170e65,
        64'h85930000_45970b50,
        64'h0613a025_04f71063,
        64'h4789873e_27810ff7,
        64'hf7932781_87aae03f,
        64'hf0ef853e_0fe00593,
        64'h43dcfd84_37830607,
        64'hb823fd84_3783d7f8,
        64'h4719fd84_37830607,
        64'ha223fd84_378302e7,
        64'h8023fd84_37830207,
        64'hc703fd04_3783cfd8,
        64'hfd843783_4fd8fd04,
        64'h3783cf98_fd843783,
        64'h4f98fd04_3783cbd8,
        64'hfd843783_4bd8fd04,
        64'h3783cb98_fd843783,
        64'h4b98fd04_3783c7d8,
        64'hfd843783_47d8fd04,
        64'h3783d3d8_1117071b,
        64'h11111737_fd843783,
        64'hc798fd84_37834798,
        64'hfd043783_c3d8fcc4,
        64'h2703fd84_378300e7,
        64'h9023fd84_37830007,
        64'hd703fd04_37831207,
        64'ha9230000_4797a62d,
        64'h478514e7_a0234705,
        64'h00004797_c61ff0ef,
        64'h1d050513_00004517,
        64'h1d058593_00004597,
        64'h0b400613_a025c7fd,
        64'hfd043783_1607a423,
        64'h00004797_cb89fd84,
        64'h3783fcf4_262387b2,
        64'hfcb43823_fca43c23,
        64'h0080f822_fc067139,
        64'h80826105_644260e2,
        64'h0001e8df_f0ef853e,
        64'h85bafea4_47039381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef40523_87bafef4,
        64'h05a387b6_fef42623,
        64'h873286ae_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e2853e,
        64'h87aae7ff_f0ef853e,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_05a387ba,
        64'hfef42623_872e87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h0001f39f_f0ef853e,
        64'h85bafe84_57039381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef41423_87bafef4,
        64'h05a387b6_fef42623,
        64'h873286ae_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e2853e,
        64'h87aaf1df_f0ef853e,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_05a387ba,
        64'hfef42623_872e87aa,
        64'h1000e822_ec061101,
        64'h80826145_74220001,
        64'hc398fd44_2703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_2a2387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61457422,
        64'h000100e7_9023fd64,
        64'h5703fe84_3783fef4,
        64'h3423fd84_3783fcf4,
        64'h1b2387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61457422_000100e7,
        64'h8023fd74_4703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_0ba387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61056462,
        64'h853e2781_439cfe84,
        64'h3783fea4_34231000,
        64'hec221101_80826105,
        64'h6462853e_93c117c2,
        64'h0007d783_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61056462,
        64'h853e0ff7_f7930007,
        64'hc783fe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826145_7422853e,
        64'hfe843783_fae7f5e3,
        64'h47850007_871bfe44,
        64'h2783fef4_22232785,
        64'hfe442783_a829fef4,
        64'h342397ba_f0c70713,
        64'h00004717_078a97ba,
        64'h078e87ba_fe446703,
        64'h02f71063_27812701,
        64'hfde45703_0007d783,
        64'h97baf3e6_8713078a,
        64'h97ba078e_87bafe44,
        64'h67030000_4697a0b9,
        64'hfe042223_fe043423,
        64'hfcf41f23_87aa1800,
        64'hf4227179_8082fea7,
        64'heee3ff87_37830200,
        64'hc737953a_02f50533,
        64'h47d1ff87_b7030200,
        64'hc7b78082_ff87b503,
        64'h0200c7b7_80826125,
        64'h70a2a1bf_f0efe43a,
        64'hecc6e8c2_e4bef406,
        64'h72c50513_567d080c,
        64'h86b21838_ec2ee0ba,
        64'hfc36ffff_f517e82a,
        64'h711da43f_f06f72e5,
        64'h0513ffff_f51785aa,
        64'h862e86b2_87368082,
        64'h610560e2_a5dff0ef,
        64'hec06a645_0513002c,
        64'h567d872e_00000517,
        64'h86aa1101_80826161,
        64'h60e2a7bf_f0efe43a,
        64'he4c6e0c2_fc3eec06,
        64'h10387745_0513f83a,
        64'hfffff517_85aa862e,
        64'h86b2f436_715d8082,
        64'h616160e2_aa5ff0ef,
        64'he43ae4c6_e0c2fc3e,
        64'hec067a25_05131018,
        64'h567df83a_f032ffff,
        64'hf51785aa_86aef436,
        64'h715d8082_612560e2,
        64'had1ff0ef_e43aecc6,
        64'he8c2e4be_ec06ae65,
        64'h0513567d_1038858a,
        64'he0baf832_f42e0000,
        64'h051786aa_fc36711d,
        64'hb31d4809_b32d4821,
        64'hbb1d4841_0206e693,
        64'hbb498da2_99020250,
        64'h051385d2_866e86ce,
        64'h001d8413_b7d58622,
        64'h2c859902_00160413,
        64'h02000513_85d286ce,
        64'hbb6d8db2_8aea018c,
        64'he563c019_fc089de3,
        64'hfff8869b_fe0a82e3,
        64'hc51901b7_06330007,
        64'h450378a2_77029902,
        64'h85d286ce_f83af03a,
        64'hf4460705_88b6b7e1,
        64'h78c28df2_8cc27762,
        64'h7e027822_99020200,
        64'h051385d2_86ce866e,
        64'hf072f442_f846fc3a,
        64'h001d8e13_b7c90785,
        64'ha08140ed_8db38cc2,
        64'h018ce863_001c881b,
        64'he4110006_841b8a89,
        64'h00060c9b_8666011c,
        64'hf3638646_000a8863,
        64'h40e78cbb_2a814006,
        64'hfa9302f6_1b63c199,
        64'h0007c583_87ba00f7,
        64'h06339381_02089793,
        64'h00088563_57fd000a,
        64'hb703008a_8d13b7cd,
        64'h8ca22b05_99020200,
        64'h051385d2_86ce001c,
        64'h84138666_b5598de6,
        64'h8aea018b_6563c019,
        64'h9902001d_8c93008a,
        64'h8d1385d2_866e86ce,
        64'h000ac503_ff8764e3,
        64'h001d8d13_00170b1b,
        64'h8dea875a_99020200,
        64'h051385d2_86ce866e,
        64'ha8094705_e00d4b05,
        64'h0006841b_8a89b7ed,
        64'h8f7d67e2_dbe50807,
        64'hf793b769_93014781,
        64'he062e436_17020ff7,
        64'h7713ca09_000aa703,
        64'h0407f613_b755e062,
        64'he4364781_000ab703,
        64'hc7191007_f713bde5,
        64'h4781e062_e436000a,
        64'hb703c719_bff1000a,
        64'ha783b7cd_000a9783,
        64'hc7810807_f793bfd9,
        64'h40e6073b_93fde062,
        64'he43600e7_c63341f7,
        64'hd71b000a_c783cf09,
        64'h0406f713_b789bb7f,
        64'hf0ef854a_85d2866e,
        64'h86ce93fd_40e60733,
        64'h00f74633_43f7d713,
        64'he062e436_000ab783,
        64'hc31d87b6_1006f713,
        64'hb5dd0780_0793eef5,
        64'h09e30750_0793a89d,
        64'h4841e03e_e436008a,
        64'h8413000a_b70347c1,
        64'h0216e693_d4f51ae3,
        64'h07000793_f0f50ce3,
        64'h06f00793_02a7e563,
        64'h12f50f63_07300793,
        64'hb71d0640_07930ef5,
        64'h06630630_0793bddd,
        64'h0c06e693_8082614d,
        64'h6da66d46_6ce67c06,
        64'h7ba67b46_7ae66a0a,
        64'h69aa694a_64ea000d,
        64'h851b740a_70aa9902,
        64'h450185d2_86cefff9,
        64'h8613013d_e463866e,
        64'hda0517e3_0004c503,
        64'h8aa28daa_cf5ff0ef,
        64'h854a85d2_866e86ce,
        64'h93fd40e6_073300f7,
        64'h463343f7_d713e062,
        64'he436000a_b783cf45,
        64'h10c51c63_06400613,
        64'h00c50663_008a8413,
        64'h02085813_270187b6,
        64'h06900613_18022006,
        64'hf7139af9_c3914006,
        64'hf7939acd_00f50363,
        64'h06400793_00f50763,
        64'h48299abd_06900793,
        64'h2ef50463_06200793,
        64'h2ef50663_06f00793,
        64'h2ef50663_05800793,
        64'h2ef50c63_07800793,
        64'he4f514e3_05800793,
        64'h2ef50863_02500793,
        64'h0ca7ef63_00f50c63,
        64'h06200793_0ea7ec63,
        64'h02f50263_00170493,
        64'h06900793_00074503,
        64'h0806e693_0ef60e63,
        64'h0014c603_a0390024,
        64'h87133006_e693a821,
        64'h1006e693_00f60563,
        64'h0014c603_b7e907a0,
        64'h061300c7_89630740,
        64'h0613bf65_84babf75,
        64'h8abe0489_28814881,
        64'h0008d363_008a8793,
        64'h000aa883_00f61d63,
        64'h02a00793_a8998726,
        64'h04c78063_06a00613,
        64'h04c78c63_06800613,
        64'h02f66d63_04c78663,
        64'h00148713_06c00613,
        64'h0004c783_fef671e3,
        64'h0ff7f793_fd07079b,
        64'h00148593_0004c703,
        64'h00e888bb_fd08889b,
        64'h84ae031b_88bbb775,
        64'h84b28aba_40f00c3b,
        64'h0026e693_0007d663,
        64'h00078c1b_008a8713,
        64'h000aa783_fce796e3,
        64'h4c0102a0_0713a825,
        64'h462584ba_06f5ee63,
        64'h4006e693_0ff7f793,
        64'hfd06079b_00148713,
        64'h45a50014_c60306f7,
        64'h17634881_02e00793,
        64'h0004c703_fef671e3,
        64'h0ff7f793_fd07079b,
        64'h00148593_0004c703,
        64'h00e30c3b_fd03031b,
        64'h84ae038b_833bbf75,
        64'h0106e693_b7c90086,
        64'he693b7e1_0046e693,
        64'hb7f90026_e693a025,
        64'h46254c01_06e5e963,
        64'h45a50ff7_7713fd07,
        64'h871b02a7_856302b7,
        64'h8463fcf7_6fe302e7,
        64'h85630014_86130004,
        64'hc78384b2_0016e693,
        64'h02879163_03000413,
        64'h02878f63_02d00413,
        64'ha8210230_05130200,
        64'h059302b0_07134681,
        64'ha15585d2_866e86ce,
        64'h001d8413_00f50863,
        64'h04850250_0793ac81,
        64'h4ba9ec3e_4d81fffb,
        64'h07936b41_cc890913,
        64'h00000917_e589892a,
        64'h8aba84b6_89b28a2e,
        64'he4eee8ea_ece6f0e2,
        64'hf4def8da_f122f506,
        64'hfcd6e152_e54ee94a,
        64'hed267171_808298df,
        64'hf06fc119_b7e1006e,
        64'h033b8082_616160a6,
        64'hd17ff0ef_887e1018,
        64'h0008089b_e43ae876,
        64'he0464746_fc579de3,
        64'hc319fe6f_0fa39f3e,
        64'h0ff37313_02010f13,
        64'h07850307_57330303,
        64'h031b03e3_ee630fff,
        64'h73130307_7f330200,
        64'h0293ff63_0e1b43a5,
        64'h47810410_0313000e,
        64'h04630610_0313020e,
        64'hfe13c721_47810003,
        64'h0463400e_f313fefe,
        64'hfe93e319_4ee68fbe,
        64'he486715d_b7e1006e,
        64'h033b8082_616160a6,
        64'hd97ff0ef_887e1018,
        64'h0008089b_e43ae876,
        64'he0464746_fc579de3,
        64'hc319fe6f_0fa39f3e,
        64'h0ff37313_02010f13,
        64'h07850307_57330303,
        64'h031b03e3_ee630fff,
        64'h73130307_7f330200,
        64'h0293ff63_0e1b43a5,
        64'h47810410_0313000e,
        64'h04630610_0313020e,
        64'hfe13c721_47810003,
        64'h0463400e_f313fefe,
        64'hfe93e319_4ee68fbe,
        64'he486715d_b7a98622,
        64'h9b020016_04130200,
        64'h051385de_86e2b791,
        64'h9b0285de_86e20009,
        64'h4503b7ed_41540cb3,
        64'h02095913_02099913,
        64'hbf89ff27_e3e3009c,
        64'h87b384ea_00148d13,
        64'h67229b02_e43a0200,
        64'h051385de_86e28626,
        64'hb7ad00d6_00230087,
        64'h0633da3d_0087f613,
        64'hbf9d02b0_06130087,
        64'h06b3c611_0047f613,
        64'hbfa10620_06130087,
        64'h06b3f886_ece346fd,
        64'hf6d898e3_4689b7bd,
        64'h05800613_008706b3,
        64'hfa86e7e3_46fd8082,
        64'h61658532_6d426ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_0b37e163,
        64'h415607b3_0209d993,
        64'h1982000a_09630094,
        64'h06330b2c_9663197d,
        64'h412d0633_01248d33,
        64'hfff70c93_00870933,
        64'hcbcd84d6_8b8d0405,
        64'h00c68023_02d00613,
        64'h008706b3_08080463,
        64'h00d40b63_02000693,
        64'h040500c6_80230300,
        64'h06130087_06b30286,
        64'he66346fd_040500c6,
        64'h80230780_06130087,
        64'h06b30486_e06346fd,
        64'head10207_f6930ad8,
        64'h966346c1_4401bf55,
        64'hfe6e0fa3_00870e33,
        64'h0405a0e9_02c89a63,
        64'h84364609_02c88163,
        64'h14794641_c285fff4,
        64'h06930286_95639281,
        64'h02099693_00868763,
        64'h92811682_cc0dee15,
        64'h4007f613_ca3d0107,
        64'hf61302b4_1e6300a4,
        64'h7463c609_03000313,
        64'h02000593_91010209,
        64'h9513fea4_69e3fe6e,
        64'h0fa30087_0e330405,
        64'h00b40963_a8010300,
        64'h03130200_05939101,
        64'h02069513_39fdc191,
        64'h00c7f593_00081563,
        64'hc6190009_89630017,
        64'hf613040a_1a6359e6,
        64'h56c68ab2_8bae8b2a,
        64'h8c362a01_e86aec66,
        64'he8caeca6_f486f062,
        64'hf45ef85a_fc560027,
        64'hfa13e4ce_e0d2478a,
        64'h843ef0a2_71598082,
        64'h8302658c_0005b303,
        64'hc5098082_808200a5,
        64'h802395b2_00d67563,
        64'hbbe102f0_00efd7e5,
        64'h05130000_6517bd35,
        64'hb4250513_85a60000,
        64'h65170470_00efb365,
        64'h05130000_6517cd09,
        64'h84aada9f_f0ef8552,
        64'h865a020a_a5830630,
        64'h00efd9a5_05130000,
        64'h6517f579_90e30804,
        64'h84930770_00ef2985,
        64'ha8850513_00006517,
        64'hff2c17e3_089000ef,
        64'h0905d3a5_05130000,
        64'h65170009_45830704,
        64'h8c130284_89130a30,
        64'h00efdc25_05130000,
        64'h65170af0_00efdb65,
        64'h05130000_6517708c,
        64'h0bd000ef_dac50513,
        64'h00006517_6c8c0cb0,
        64'h00efda25_05130000,
        64'h6517688c_ff2c17e3,
        64'h0dd000ef_0905d8e5,
        64'h05130000_65170009,
        64'h45830109_0c130f30,
        64'h00efdaa5_05130000,
        64'h6517fe99_17e31030,
        64'h00ef0905_db450513,
        64'h00006517_00094583,
        64'hff048913_119000ef,
        64'hda850513_00006517,
        64'h125000ef_d9e50513,
        64'h85ce0000_6517bf15,
        64'hd8a50513_85ce0000,
        64'h651713f0_00efc2e5,
        64'h05130000_6517cd09,
        64'h4b910804_89aa8a8a,
        64'hea7ff0ef_850a4605,
        64'h710144ac_161000ef,
        64'hd9850513_00006517,
        64'h45d616f0_00efd865,
        64'h05130000_651745c6,
        64'h17d000ef_d6c50513,
        64'h00006517_65a618b0,
        64'h00efd625_05130000,
        64'h65177582_199000ef,
        64'hd5850513_00006517,
        64'h65e21a70_00efd4e5,
        64'h05130000_651745d2,
        64'h1b5000ef_d4450513,
        64'h00006517_45c21c30,
        64'h00efd3a5_05130000,
        64'h651745b2_1d1000ef,
        64'hd3050513_00006517,
        64'h45a21df0_00efd265,
        64'h05130000_65176582,
        64'h1ed000ef_d1450513,
        64'h00006517_b75554f9,
        64'h1fd000ef_d0450513,
        64'h00006517_fa843583,
        64'h20d000ef_cfc50513,
        64'h00006517_faa43423,
        64'hc11df71f_f0ef848a,
        64'h850a4585_46057101,
        64'h22d000ef_d0450513,
        64'h00006517_80826125,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h64468526_60e6fa04,
        64'h011354fd_259000ef,
        64'hd0850513_00006517,
        64'hc51df39f_f0ef8b2e,
        64'h8a2a1080_e862ec5e,
        64'hf456fc4e_e0cae4a6,
        64'hec86f05a_f852e8a2,
        64'h711d8082_014160a2,
        64'h557d28f0_00efd1e5,
        64'h05130000_651785aa,
        64'hc90921d0_20efe406,
        64'hc0c50513_46051141,
        64'h00005517_86aab76d,
        64'h45012b70_00efd265,
        64'h05130000_6517bf6d,
        64'h55752c70_00efd065,
        64'h05130000_6517c909,
        64'h85aa71c0_10ef8522,
        64'hbfd15579_2e1000ef,
        64'hcf850513_00006517,
        64'hc90985aa_651000ef,
        64'h852285aa_c5c40413,
        64'h00005417_41508082,
        64'h01416402_60a2557d,
        64'h30d000ef_d0450513,
        64'h00006517_ed014270,
        64'h00ef4501_321000ef,
        64'he022e406_d0650513,
        64'h11410000_65178082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_00a78223,
        64'h0ff57513_00d78023,
        64'h0085551b_0ff57693,
        64'h00d78623_f8000693,
        64'h00078223_01e71793,
        64'h470d02b5_553b0045,
        64'h959b8082_00a78023,
        64'hdf650207_77130147,
        64'hc70307fa_478d8082,
        64'h02057513_0147c503,
        64'h07fa478d_80820005,
        64'h45038082_00b50023,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_100004b7,
        64'h1c858593_00005597,
        64'hf1402573_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_415040ef,
        64'h40000137_03249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
