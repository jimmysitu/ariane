/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 2107;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00000078_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000078_36313025,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000078_36313025,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_78323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000a64_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h00000a64_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_0000000a,
        64'h78363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h0000000a_78363130,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h0000000a_78363130,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_00000a64,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_00000a64,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_00000a64,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_00000a64,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h00000000_00000a78,
        64'h25202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h00000000_0a642520,
        64'h3a737574_61747320,
        64'h2c64656c_69616620,
        64'h64616552_20304453,
        64'h00000000_0a216465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a6425,
        64'h203a7375_74617473,
        64'h202c6465_6c696166,
        64'h206e6f69_74617a69,
        64'h6c616974_696e6920,
        64'h64726163_20304453,
        64'h0000000a_6425203a,
        64'h73757461_7473202c,
        64'h64656c69_6166206c,
        64'h61697469_6e692067,
        64'h69666e6f_63204453,
        64'h00000000_0000000a,
        64'h2164656c_69616620,
        64'h6769666e_6f632070,
        64'h756b6f6f_6c204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_002e2e2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd0080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h08090000_38000000,
        64'hda0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000a001,
        64'h824fe0ef_19c50513,
        64'h00001517_84025965,
        64'h85930000_05971000,
        64'h0437e901_dbefd0ef,
        64'h10000537_65a184af,
        64'he0ef21a5_05130000,
        64'h1517856f_e0ef1c65,
        64'h05130000_1517950f,
        64'he0ef2404_051386af,
        64'he0ef1da5_05130000,
        64'h1517964f_e0ef2404,
        64'h0513000f_4437882f,
        64'he0ef1ca5_05130000,
        64'h1517d1cf_d0efe022,
        64'he406a005_05132005,
        64'h85931141_02626537,
        64'h65f18082_0141421c,
        64'h920100f6_90231602,
        64'h47892641_640260a2,
        64'h80820141_45056402,
        64'h60a28082_01414505,
        64'h00f61023_3ff7879b,
        64'h920177fd_16026402,
        64'h60a20326_061bfe07,
        64'h56e38b89_4107571b,
        64'h0107971b_93c117c2,
        64'h0006d783_ef9da011,
        64'h92811682_0306069b,
        64'h4050e129_de0fe0ef,
        64'h842ae406_e0226000,
        64'h05934681_862e1141,
        64'h80820141_439c9381,
        64'h00e69023_17824709,
        64'h0106079b_640260a2,
        64'h80820141_450562e7,
        64'ha2234705_00000797,
        64'h640260a2_948fe0ef,
        64'h67050513_68458593,
        64'h35c00613_00001517,
        64'h00001597_80820141,
        64'h45056402_60a28082,
        64'h01414505_64e7ad23,
        64'h47050000_07976402,
        64'h60a297ef_e0ef6a65,
        64'h05136ba5_859335d0,
        64'h06130000_15170000,
        64'h15978082_01414505,
        64'h00e79023_3ff7071b,
        64'h9381777d_17826402,
        64'h60a20326_079bfe07,
        64'h56e38b89_4107571b,
        64'h0107971b_93c117c2,
        64'h0006d783_ebd9a011,
        64'h92811682_0306069b,
        64'h4050e53d_eb0fe0ef,
        64'h6ce79a23_85228005,
        64'h85934601_46854745,
        64'h00000797_6585c0df,
        64'he0ef8522_458500e7,
        64'h90239381_17822791,
        64'h862e2000_0713405c,
        64'hfee79de3_07850007,
        64'h802308d6_12632005,
        64'h871387ae_842a1116,
        64'h86937007_a9231111,
        64'h16b70000_07975150,
        64'hc979e022_e4061141,
        64'h80820141_853e4785,
        64'h72e7a723_47050000,
        64'h07976402_60a2a52f,
        64'he0ef77a5_051378e5,
        64'h859332c0_06130000,
        64'h15170000_15978082,
        64'h0141853e_00a037b3,
        64'h640260a2_f50fe0ef,
        64'ha0058593_46014681,
        64'h852265ad_f17d4785,
        64'hf64fe0ef_70058593,
        64'h4681658d_49308082,
        64'h0141853e_640260a2,
        64'h478578e7_a8234705,
        64'h00000797_ab0fe0ef,
        64'h7d850513_7ec58593,
        64'h32d00613_00001517,
        64'h00001597_02f70963,
        64'h842a1117_87931111,
        64'h17b77c07_a0235158,
        64'h00000797_cd25e022,
        64'he4061141_bd85bd8f,
        64'he0ef4505_dc0780e3,
        64'h0807f793_0007d783,
        64'hb3f14505_7ee7a523,
        64'h47050000_0797b0af,
        64'he0ef8325_05138465,
        64'h859348e0_06130000,
        64'h25170000_2597b7e9,
        64'hffcfe0ef_85d2fd37,
        64'h98e38522_85ca4601,
        64'h46850344_4783c0a1,
        64'hc3290407_77130007,
        64'hd7039381_178203e7,
        64'h879b405c_e20510e3,
        64'h0ff4f493_34fd833f,
        64'he0efa01d_300a0a13,
        64'h4985c54f_e0ef00e7,
        64'h90230407_67130280,
        64'h0493500a_09130007,
        64'hd7039381_86d71723,
        64'h46c10000_17171782,
        64'h00d71023_03e7879b,
        64'h93011702_0047871b,
        64'h45056a05_405c0400,
        64'h069300f7_04630800,
        64'h0693478d_03744703,
        64'h08f71b63_11178793,
        64'h111117b7_8a07a523,
        64'h50580000_1797bd69,
        64'h4505d939_c63ff0ef,
        64'h85225005_8593dc1c,
        64'h031975b7_5007879b,
        64'h031977b7_00f69023,
        64'h4789bd7d_4505dd2d,
        64'hc87ff0ef_85220805,
        64'h8593dc1c_02faf5b7,
        64'h0807879b_02faf7b7,
        64'h00f69023_4789b5a5,
        64'hfe0756e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d783ef9d,
        64'ha0119281_16820306,
        64'h069b4050_f00514e3,
        64'h915fe0ef_60000593,
        64'h10060613_468103b9,
        64'h0637b5f5_439c9381,
        64'h178227c1_405c00e7,
        64'h80230047_67130007,
        64'hc7039381_17820287,
        64'h879b4501_405cd60f,
        64'he0ef3e80_05130af7,
        64'h0a63479d_5478f921,
        64'hd17ff0ef_852200f6,
        64'h90234789_5c0cb5e5,
        64'hfe0756e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d783efc9,
        64'ha0119281_16820306,
        64'h069b4050_f159993f,
        64'he0ef9ae7_9b238522,
        64'h60000593_16454685,
        64'h47450000_17978100,
        64'h0637ef1f_e0ef4585,
        64'h00e79023_93811782,
        64'h2791860a_04000713,
        64'h415c8082_61654505,
        64'h6a0669a6_694664e6,
        64'h9ee7a323_47050000,
        64'h17977406_70a6d0af,
        64'he0efa325_0513a465,
        64'h85931f30_06130000,
        64'h25170000_25978082,
        64'h61656a06_69a66946,
        64'h64e67406_70a64505,
        64'hd135a0ff_e0ef8522,
        64'h60000593_46812006,
        64'h0613dd1c_03b90637,
        64'h2007879b_0bebc7b7,
        64'h80826165_6a0669a6,
        64'h694664e6_740670a6,
        64'h4505a4e7_a8234705,
        64'h00001797_d70fe0ef,
        64'ha9850513_aac58593,
        64'h1f400613_00002517,
        64'h00002597_80826165,
        64'h45056a06_69a66946,
        64'h64e600f6_10233ff7,
        64'h879b9201_77fd1602,
        64'h740670a6_0326061b,
        64'hfe0755e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d7831207,
        64'h9a63a019_92811682,
        64'h0306069b_4050e145,
        64'haadfe0ef_85226000,
        64'h05934681_10060613,
        64'hdd1c03b9_06375007,
        64'h879b0319_77b70af7,
        64'h0163479d_55781ae7,
        64'h88634709_10e78b63,
        64'h47050345_478308f7,
        64'h1363842a_11178793,
        64'h111117b7_b007a123,
        64'h51580000_17971005,
        64'h0263fc02_f802f402,
        64'hf002ec02_e802e402,
        64'he002e0d2_e4cee8ca,
        64'heca6f0a2_f4867159,
        64'h80820141_4505b2e7,
        64'haa234705_00001797,
        64'h60a2e56f_e0efb7e5,
        64'h0513b925_85932b70,
        64'h06130000_25170000,
        64'h2597b75d_00c69023,
        64'h92411642_8e5d0622,
        64'h8fd90017_e7938205,
        64'h03f7f793_071a0096,
        64'h57130006_d783fee5,
        64'he8e32785_92410307,
        64'h961302f8_573bf8a7,
        64'h8be3a019_7ff00513,
        64'h47858082_014100f6,
        64'h90230047_e7934501,
        64'h60a20006_d783dfed,
        64'h8b890006_d78300e6,
        64'h90239341_17428f5d,
        64'h0017e793_0ff7f793,
        64'h07228305_0006d783,
        64'hbfd9bce7_a8234705,
        64'h00001797_ef0fe0ef,
        64'hc1850513_c2c58593,
        64'h2b800613_00002517,
        64'h00002597_80820141,
        64'h450560a2_f6759341,
        64'h03051713_02f5fc63,
        64'h367d0017_151b02e8,
        64'h57bb0717_8e630365,
        64'h478300f6_902393c1,
        64'h17c29be9_93c117c2,
        64'h47054625_0006d783,
        64'h92811682_02c6869b,
        64'h48890085_28034154,
        64'h04f71863_11178793,
        64'h111117b7_c407a523,
        64'h51580000_17971005,
        64'h0063e406_11418082,
        64'h0141439c_938100e6,
        64'h90231782_47090106,
        64'h079b6402_60a28082,
        64'h01414505_c6e7ad23,
        64'h47050000_17976402,
        64'h60a2f9ef_e0efcc65,
        64'h0513cda5_859319f0,
        64'h06130000_25170000,
        64'h25978082_01414505,
        64'h640260a2_80820141,
        64'h4505cae7_a8234705,
        64'h00001797_640260a2,
        64'hfd4fe0ef_cfc50513,
        64'hd1058593_1a000613,
        64'h00002517_00002597,
        64'h80820141_450500e7,
        64'h90233ff7_071b9381,
        64'h777d1782_640260a2,
        64'h0326079b_fe0756e3,
        64'h8b894107_571b0107,
        64'h971b93c1_17c20006,
        64'hd783ebd9_a0119281,
        64'h16820306_069b4050,
        64'he53dd07f_e0efd2e7,
        64'h95238522_60000593,
        64'h16414685_47450000,
        64'h17970100_0637a64f,
        64'hf0ef8522_458500e7,
        64'h90239381_17822791,
        64'h862e0400_0713405c,
        64'hfee79de3_07850007,
        64'h802308d6_13630405,
        64'h871387ae_842a1116,
        64'h8693d607_a5231111,
        64'h16b70000_17975150,
        64'hcd61e022_e4061141,
        64'hb76500e6_90230047,
        64'h67139b61_93411742,
        64'h0006d703_92811682,
        64'h03e7869b_405cb5fd,
        64'h4505d551_d91fe0ef,
        64'h85226005_85934609,
        64'h468102f4_0ba365a1,
        64'h4789f005_15e3dabf,
        64'he0ef8522_70058593,
        64'h4681658d_4830b7a9,
        64'h4501439c_93811782,
        64'h27c1405c_04f70163,
        64'h47915478_00e78023,
        64'h0ff77713_0206e713,
        64'h00c59463_0026e713,
        64'h0ff6f693_0007c683,
        64'h93811782_0287879b,
        64'h460d0374_4583405c,
        64'ha13fe0ef_3e800513,
        64'h00f69023_4789b725,
        64'h60078613_f2e698e3,
        64'h20078613_471102e4,
        64'h0ba303b7_07b7470d,
        64'hf2f718e3_47a14858,
        64'h80820141_4505e4e7,
        64'ha2234705_00001797,
        64'h640260a2_969fe0ef,
        64'he9050513_ea458593,
        64'h11200613_00002517,
        64'h00002597_b7e5f4e7,
        64'he1e34501_478d4958,
        64'hb7495007_86138082,
        64'h01416402_60a24505,
        64'he8e7a323_47050000,
        64'h17979a7f_e0efece5,
        64'h0513ee25_85931130,
        64'h06130000_25170000,
        64'h25978082_01416402,
        64'h60a24505_00f61023,
        64'h3ff7879b_920177fd,
        64'h16020326_061bfe07,
        64'h56e38b89_4107571b,
        64'h0107971b_93c117c2,
        64'h0006d783_e3e1a011,
        64'h92811682_0306069b,
        64'h4050ed05_ed9fe0ef,
        64'h85226000_05934681,
        64'h06e68f63_10078613,
        64'h471102e4_0ba303b7,
        64'h07b74709_0ce78863,
        64'h54740752_20005737,
        64'h8ff91782_0ff78793,
        64'h00ff07b7_781814f7,
        64'h0e634785_03444703,
        64'h0af70e63_47890365,
        64'h470308f7_1a63842a,
        64'h11178793_111117b7,
        64'hf407a323_51580000,
        64'h1797c565_e022e406,
        64'h1141b7a9_439c9381,
        64'h00e69023_17824709,
        64'h0106079b_80826105,
        64'h450564a2_f6e7a923,
        64'h47050000_17976442,
        64'h60e2a97f_e0effbe5,
        64'h0513fd25_85930b90,
        64'h06130000_25170000,
        64'h2597bfb1_450500e7,
        64'h90233ff7_071b9381,
        64'h777d1782_0326079b,
        64'hfe0756e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d783efb1,
        64'ha0119281_16820306,
        64'h069b4050_f951fc3f,
        64'he0effee7_93238522,
        64'h30058593_46014685,
        64'h47450000_179765ad,
        64'hd1eff0ef_85224585,
        64'h00e79023_93811782,
        64'h27918626_4721405c,
        64'h80826105_64a26442,
        64'h60e24505_00e7a923,
        64'h47050000_1797b33f,
        64'he0ef05a5_051306e5,
        64'h85930ba0_06130000,
        64'h25170000_25978082,
        64'h610564a2_644260e2,
        64'h4505cd15_830ff0ef,
        64'h85227005_85934681,
        64'h658d4830_fee79de3,
        64'h07850007_802302d6,
        64'h16630085_871387ae,
        64'h84ae842a_11168693,
        64'h0607a823_111116b7,
        64'h00001797_5150c17d,
        64'he426e822_ec061101,
        64'h80826105_450564a2,
        64'h08e7a723_47050000,
        64'h17976442_60e2bb3f,
        64'he0ef0da5_05130ee5,
        64'h859307e0_06130000,
        64'h25170000_2597b765,
        64'h00979023_43189381,
        64'h8cf59301_17821702,
        64'h27910107_871b16fd,
        64'h6685405c_f1718c2f,
        64'hf0ef6585_4681862e,
        64'h84aebfc9_0ee7a123,
        64'h47050000_1797c03f,
        64'he0ef12a5_051313e5,
        64'h859307f0_06130000,
        64'h25170000_25978082,
        64'h610564a2_644260e2,
        64'h4505cb8d_3037f793,
        64'h439c9381_17820247,
        64'h879b415c_02f71163,
        64'h842a1117_87931111,
        64'h17b71207_a8235158,
        64'h00001797_c541e426,
        64'he822ec06_1101b6c1,
        64'h4905ea05_01e31f80,
        64'h00ef8522_b6f94905,
        64'heaf708e3_47890b94,
        64'hc703b5c1_c4079de3,
        64'h0a24c783_00e78e63,
        64'h4711bcd7_13e30b94,
        64'hc703bd39_02f40e23,
        64'h4785d85f_e0ef00e7,
        64'h90230047_67133e80,
        64'h05130007_d703b901,
        64'h4905def7_09e34785,
        64'h0b94c703_be051ce3,
        64'h285000ef_852285a6,
        64'hc00512e3_688000ef,
        64'h8522d47c_4795bfd5,
        64'h93411742_0007d703,
        64'heb158b09_93411742,
        64'h0007d703_00e79023,
        64'h00176713_0007d703,
        64'h93811782_02c7879b,
        64'hc2070ee3_8b210007,
        64'h57039301_170203e7,
        64'h871b405c_dfffe0ef,
        64'h00e79023_00876713,
        64'h0007d703_00e69023,
        64'h93819341_17429b69,
        64'h93411742_178203e7,
        64'h879b0006_d7039281,
        64'h168202c7_869b3885,
        64'h05136505_405cec07,
        64'h9ee303c4_4783eef7,
        64'h12e347a1_4858eee7,
        64'hf6e3478d_00d14703,
        64'hbfbdd47c_4795fee7,
        64'hf5e34785_03744703,
        64'hdbed8b89_bba1d3f1,
        64'h0a24c783_d47c4799,
        64'hc71900c7_f713b755,
        64'hd47c4791_00f9f863,
        64'h03744783_c30d00c7,
        64'hf713b311_892ab321,
        64'h4905ee05_05e34930,
        64'h00ef8522_10058593,
        64'h03a205b7_ee079ee3,
        64'h0a24c783_12e6fb63,
        64'h4685ffc7_871b14e7,
        64'h8c63471d_547cd005,
        64'h19e339f0_00ef8522,
        64'h85a6d005_1fe37a20,
        64'h00ef8522_d47c479d,
        64'h06e9f363_03744703,
        64'hcf210307_f7130c44,
        64'hc783d07c_8fd90d44,
        64'hc703d07c_8fd90087,
        64'h171b0d54_c703d07c,
        64'h27818fd9_0107979b,
        64'h0d64c783_d0780187,
        64'h971b0d74_c783d605,
        64'h15e33f70_00ef11c4,
        64'h84938522_11c48593,
        64'h00001497_d80510e3,
        64'h3da000ef_8522bb45,
        64'h4905d941_011000ef,
        64'h8522d47c_4795f8e7,
        64'hffe34785_03744703,
        64'hd3dd8b89_00d14783,
        64'hd7dd0004_c7831007,
        64'hc9630024_8783ed69,
        64'h5ec000ef_8522858a,
        64'hdc0512e3_41e000ef,
        64'h8522c791_8b910014,
        64'hc783dc05_1be33020,
        64'h00ef8522_85a6de05,
        64'h11e33c30_00ef8522,
        64'hbd09e8f7_08e34785,
        64'h03444703_e8f71de3,
        64'h47915478_1efa6963,
        64'h03744783_c7898b89,
        64'h0c44c783_d07c8fd9,
        64'h0d44c703_d07c8fd9,
        64'h0087171b_0d54c703,
        64'hd07c2781_8fd90107,
        64'h979b0d64_c783d078,
        64'h0187971b_0d74c783,
        64'he2051ee3_4c9000ef,
        64'h1ee48493_85221ee4,
        64'h85930000_1497e405,
        64'h19e34ac0_00ef8522,
        64'hef3a1be3_03644a03,
        64'heee7ffe3_478d0354,
        64'h4703bdd9_ac058593,
        64'hdc1c0121_f5b7ac07,
        64'h879b0121_f7b7bf85,
        64'h02f40a23_4789bdcd,
        64'h84058593_dc1c017d,
        64'h85b78407_879b017d,
        64'h87b702f7_00634789,
        64'h03644703_ea0514e3,
        64'hde6ff0ef_8522f0d7,
        64'h11e3bdf1_4905f0f7,
        64'h05e34795_00f6f763,
        64'h0ff7f793_fff7079b,
        64'h46850344_4703ffed,
        64'h8b890007_47839301,
        64'h170202f7_071b4058,
        64'h00e78023_47099381,
        64'h00d71023_17823ff6,
        64'h869b9301_76fd02f7,
        64'h879b1702_00c69023,
        64'h0327871b_92811682,
        64'h0307869b_567d405c,
        64'h02f40a23_4785c949,
        64'hcb4ff0ef_85221000,
        64'h059340ff_86374681,
        64'hbf894905_4ce7ad23,
        64'h47050000_1797ffbf,
        64'he0ef5225_051351e5,
        64'h859323f0_06130000,
        64'h25170000_2597bfa5,
        64'h00a03933_3c2000ef,
        64'h85222000_0593f8f7,
        64'h05e34791_54781ee7,
        64'h82634715_10e78363,
        64'h47091937_87634985,
        64'h03444783_fd3d892a,
        64'hd1cff0ef_85227000,
        64'h05934681_4830f941,
        64'h0e7000ef_8522a805,
        64'h8593dc1c_018cc5b7,
        64'ha807879b_018cc7b7,
        64'hf54dd55f_f0ef8522,
        64'h02f50a23_4795fae7,
        64'h91e38ff5_40000737,
        64'hc00006b7_551c8082,
        64'h610d7a46_79e6690a,
        64'h64aa854a_644a60ea,
        64'h490558e7_a4234705,
        64'h00001797_8a8ff0ef,
        64'h5d050513_5cc58593,
        64'h24000613_00002517,
        64'h00002597_a01d4905,
        64'hcd69d9ef_f0ef8522,
        64'h45814601_46819c0f,
        64'hf0ef7105_05136509,
        64'h04f70b63_47890205,
        64'h0e23dd1c_a807879b,
        64'h000627b7_03654703,
        64'h02f50a23_02f50ba3,
        64'h478504f7_1163842a,
        64'h11178793_111117b7,
        64'h5e07ab23_51580000,
        64'h17971005_0463fc02,
        64'hf802f402_f002ec02,
        64'he802e402_e0020004,
        64'hb0239881_f8d2fcce,
        64'he14ae922_ed0605f1,
        64'h0493e526_7135b5f1,
        64'hd07c02e4_0aa30097,
        64'hd79b00f6_f7130126,
        64'h569b00e7_97bb00f6,
        64'hf71300e7_97bb2785,
        64'h0086d69b_27098b1d,
        64'h8fcd4210_0077571b,
        64'h8fe59201_0167559b,
        64'h160200a6_979b2681,
        64'h270101c7_861b4294,
        64'h43184210_92819301,
        64'h92011682_17021602,
        64'h0187869b_0147871b,
        64'h0107861b_c0048493,
        64'h405cf005_15e3e8af,
        64'hf0ef8522_90048593,
        64'h46816485_4830fd11,
        64'he9cff0ef_30000593,
        64'h12340637_c83cc438,
        64'h123407b7_c47cc070,
        64'hc02c0007_d7830007,
        64'h57030006_56030005,
        64'hd5839381_93019201,
        64'h91811782_17021602,
        64'h158227f1_0187871b,
        64'h0147861b_0107859b,
        64'h85224681_405cf535,
        64'heecff0ef_85222000,
        64'h05934601_4681d81c,
        64'h47850007_54630217,
        64'h97138082_61054505,
        64'h64a272e7_a0234705,
        64'h00001797_644260e2,
        64'ha44ff0ef_76c50513,
        64'h76858593_67000613,
        64'h00002517_00002597,
        64'hb751f6e7_98e38ff5,
        64'h40000737_c00006b7,
        64'h551c8082_610564a2,
        64'h644260e2_450576e7,
        64'ha2234705_00001797,
        64'ha84ff0ef_7ac50513,
        64'h7a858593_67100613,
        64'h00002517_00002597,
        64'h80826105_450564a2,
        64'h644260e2_d165f82f,
        64'hf0ef8522_10000593,
        64'h40ff8637_46810807,
        64'hc8632781_439c9381,
        64'h178227c1_405ca015,
        64'hc911fa6f_f0ef8522,
        64'h45814601_46810207,
        64'h5b6302f7_9713439c,
        64'h93811782_0247879b,
        64'h405ccb99_445c08f7,
        64'h04634789_03654703,
        64'h06f71263_842a1117,
        64'h87931111_17b77e07,
        64'haa235158_00001797,
        64'hcd4de426_e822ec06,
        64'h11018082_61454501,
        64'h69a26942_64e200f6,
        64'h90234789_740270a2,
        64'hb775dd25_811ff0ef,
        64'h82e79a23_85228005,
        64'h8593864e_4685470d,
        64'h00002797_6589b799,
        64'hf4c713e3_01077733,
        64'h40000637_c0000837,
        64'h5518bff9_f4064fe3,
        64'h02f71613_43189301,
        64'h17020247_871b8082,
        64'h61454505_69a26942,
        64'h64e27402_70a200f6,
        64'h10233ff7_879b9201,
        64'h77fd1602_0326061b,
        64'hfe0756e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d783e3c1,
        64'ha0119281_16820306,
        64'h069b4050_ed0589bf,
        64'hf0ef8ce7_90238522,
        64'h90058593_864e86a6,
        64'h02700713_00002797,
        64'h658908f4_88634785,
        64'hdffff0ef_852285a6,
        64'h864ae13d_79a000ef,
        64'h20000593_00f70763,
        64'h842a89ae_89362000,
        64'h0713439c_93811782,
        64'h2791eb59_45580ae8,
        64'h0863415c_84b24709,
        64'h03654803_e44ee84a,
        64'hf022f406_ec267179,
        64'h80826145_4501421c,
        64'h69a26942_64e29201,
        64'h00f69023_16024789,
        64'h26417402_70a2b775,
        64'hdd25927f_f0ef94e7,
        64'h95238522_10058593,
        64'h864e4685_474d0000,
        64'h27976585_b799f4c7,
        64'h13e30107_77334000,
        64'h0637c000_08375518,
        64'hbff9f406_4fe302f7,
        64'h16134318_93011702,
        64'h0247871b_80826145,
        64'h450569a2_694264e2,
        64'h740270a2_00f61023,
        64'h3ff7879b_920177fd,
        64'h16020326_061bfe07,
        64'h56e38b89_4107571b,
        64'h0107971b_93c117c2,
        64'h0006d783_e3c1a011,
        64'h92811682_0306069b,
        64'h4050ed05_9b1ff0ef,
        64'h9ce79b23_85222005,
        64'h8593864e_86a60370,
        64'h07130000_27976585,
        64'h08f48863_4785f15f,
        64'hf0ef8522_85a6864a,
        64'he13d0b10_00ef2000,
        64'h059300f7_0763842a,
        64'h89ae8936_20000713,
        64'h439c9381_17822791,
        64'heb594558_0ae80863,
        64'h415c84b2_47090365,
        64'h4803e44e_e84af022,
        64'hf406ec26_71798082,
        64'h00a8a023_08b79123,
        64'h0208d893_0805051b,
        64'h08e79023_08c7a223,
        64'h18820230_071397aa,
        64'h0588889b_83f50206,
        64'h97930265_85bb9e39,
        64'h01e7073b_7741ff07,
        64'h18e307a1_00ee073b,
        64'h00079123_01d79023,
        64'hc3d86e41_02100e93,
        64'h873201e8_083b0805,
        64'h079300c8_083b0107,
        64'h1f1b7841_ce85fff7,
        64'h069b0016_871bc399,
        64'h0006871b_93c117c2,
        64'h0107d69b_04e86963,
        64'h0007881b_468102b3,
        64'h07bb00f3_73332601,
        64'h67410007_d7839381,
        64'h17820048_879b137d,
        64'h63050045_28838082,
        64'h014100a0_353360a2,
        64'hacdff0ef_e4067000,
        64'h05934681_11414930,
        64'hb339d07c_0097d79b,
        64'h00f717bb_00f67793,
        64'h00f7173b_0086561b,
        64'h27052789_8b9d8f55,
        64'h0077d79b_8f650167,
        64'hd69bc004_849300a6,
        64'h171bb381_d07c00a7,
        64'h979b2785_93a9178a,
        64'hd4d718e3_4685cb19,
        64'h8b0d0166_d71b2601,
        64'h0007079b_43944290,
        64'h43189301_93819281,
        64'h42101782_16821702,
        64'h920127f1_16020187,
        64'h869b0147_871b0107,
        64'h861b405c_d4051be3,
        64'hb5dff0ef_85229004,
        64'h85934681_6485b599,
        64'h02f40aa3_4789bb85,
        64'h4505d16d_b79ff0ef,
        64'h85223000_05934601,
        64'h4681ee19_c8308e65,
        64'h43909381_178227c1,
        64'h405ca809_c47cc438,
        64'hc074c030_0007d783,
        64'h00075703_0006d683,
        64'h00065603_93819301,
        64'h92819201_17821702,
        64'h16821602_27f10187,
        64'h871b0147_869b0107,
        64'h861b74c1_405cdc05,
        64'h18e3bd7f_f0ef8522,
        64'h20000593_46014681,
        64'hde0491e3_fed79ee3,
        64'h8ff1431c_00d78663,
        64'h8ff1431c_93011702,
        64'h0247071b_01f006b7,
        64'h01f00637_4058821f,
        64'hf0ef00f7_10230047,
        64'he7933e80_05130007,
        64'h5783dfed_8b890007,
        64'h578300f7_10230017,
        64'he7930007_57839301,
        64'h02079713_02c7879b,
        64'he2070de3_8b210007,
        64'h57039301_170203e7,
        64'h871b405c_867ff0ef,
        64'h00f69023_0087e793,
        64'h38850513_65050006,
        64'hd7839281_00f71023,
        64'h93c117c2_9be993c1,
        64'h17c21682_03e6869b,
        64'h00075783_93011702,
        64'h02c6871b_fff58ff1,
        64'h431cc781_8ff1431c,
        64'h93011702_0246871b,
        64'h84aa01f0_06374054,
        64'hca5ff0ef_8522b005,
        64'h85934601_468102f4,
        64'h0e236585_47850c07,
        64'h5d630277_9713d818,
        64'h47050007_54630217,
        64'h9713bf75_41ff8637,
        64'hfd4792e3_485cfd37,
        64'h95e340ff_86378522,
        64'h03644783_ee0513e3,
        64'h85a64681_cf1ff0ef,
        64'h85224601_85ca4681,
        64'h0207c963_2781439c,
        64'h93811782_27c1405c,
        64'hf00515e3_d11ff0ef,
        64'ha8299004_84934a21,
        64'h49897009_091364ad,
        64'h690d02f4_0aa34785,
        64'h1af70f63_1aa00713,
        64'h431c9301_17022741,
        64'h40588082_61454505,
        64'h6a0269a2_694264e2,
        64'hd4e7af23_47050000,
        64'h27977402_70a2883f,
        64'hf0efdaa5_0513da65,
        64'h85931610_06130000,
        64'h35170000_3597b785,
        64'hf4e796e3_8ff54000,
        64'h0737c000_06b7551c,
        64'ha0a9ffed_8b890006,
        64'hc7839281_168202f7,
        64'h069b4058_00a78023,
        64'h93811782_02f7879b,
        64'h405cfaf5_12e34789,
        64'hc925daff_f0ef8522,
        64'h80058593_1aa00613,
        64'h46816585_80826145,
        64'h6a0269a2_694264e2,
        64'h740270a2_4505dee7,
        64'ha2234705_00002797,
        64'h905ff0ef_e2c50513,
        64'he2858593_16200613,
        64'h00003517_00003597,
        64'h80826145_6a0269a2,
        64'h694264e2_740270a2,
        64'h4505c521_e09ff0ef,
        64'h85224581_46014681,
        64'h00075963_02f79713,
        64'h439c9381_17820247,
        64'h879b405c_cb99445c,
        64'h0af70663_4789c95c,
        64'h47910365_470304f7,
        64'h1563842a_11178793,
        64'h111117b7_e407ad23,
        64'h51580000_2797c16d,
        64'he052e44e_e84aec26,
        64'hf022f406_7179b769,
        64'h00e79023_25013ff7,
        64'h071b777d_4509e311,
        64'hffe57713_91411542,
        64'h0007d503_93810205,
        64'h17930325_051b8082,
        64'h61054505_690264a2,
        64'heae7a323_47050000,
        64'h27976442_60e29cbf,
        64'hf0efef25_0513eee5,
        64'h859344b0_06130000,
        64'h35170000_3597b76d,
        64'h00f61023_02000793,
        64'hd6dd0206_f6930006,
        64'h56838082_61056902,
        64'h64a26442_60e24505,
        64'heee7a723_47050000,
        64'h2797a0ff_f0eff365,
        64'h0513f325_859344c0,
        64'h06130000_35170000,
        64'h35978082_61054501,
        64'h690264a2_00f61023,
        64'h47856442_60e2d7e5,
        64'h0805c763_c7318b85,
        64'h4105d59b_0107959b,
        64'h93c117c2_00065783,
        64'h92011602_0305061b,
        64'h40c800a9_20230209,
        64'h59138d5d_19028d75,
        64'h29313fff_06b70105,
        64'h151bf627_d7830000,
        64'h2797efb5_02057793,
        64'hc7818b89_439c9381,
        64'h17820249_079bcb19,
        64'h25012701_dff77713,
        64'h9f21d007_071b777d,
        64'he0bff0ef_00e79023,
        64'h93813ff7_071b777d,
        64'h178200d7_10230329,
        64'h079b9301_17020309,
        64'h071b0045_2903c390,
        64'h93811782_27a1842e,
        64'h56fd415c_00e78023,
        64'h47399381_00d71023,
        64'h17829301_92c102e7,
        64'h879b1702_16c20067,
        64'h871beb75_8b054318,
        64'h93011702_0247871b,
        64'h415c0ef7_126384aa,
        64'h11178793_111117b7,
        64'hfe07af23_51580000,
        64'h27971405_0063e04a,
        64'he426e822_ec061101,
        64'h8082bdf9_852ef4f5,
        64'h85e3c007_8793f8e5,
        64'h8de31007_8713f4f5,
        64'h8de38082_83a78513,
        64'heee68fe3_81a78513,
        64'h47050345_46838082,
        64'h31b00513_808261b0,
        64'h0513f0f7_0ce363a0,
        64'h05134785_03454703,
        64'hb715852e_fcf58ce3,
        64'h80078793_f8d58ce3,
        64'h40068693_fee584e3,
        64'h90078713_6789feb7,
        64'h71e3fee5_8be37007,
        64'h87138082_03a5e513,
        64'hf4f59ae3_50078793,
        64'h00e58663_30078713,
        64'hb78dfce5_87e3d007,
        64'h0713f6f5_88e361a5,
        64'h05136005_07936521,
        64'h8082f6f5_9fe32090,
        64'h05132000_0793f8f5,
        64'h86e31020_05131000,
        64'h07938082_01a5e513,
        64'hf8f59ee3_a0078793,
        64'hfae583e3_90978513,
        64'h90078713_0ab76f63,
        64'h00e58e63_b0078713,
        64'h8082fae5_9fe39027,
        64'h85139007_8713fce5,
        64'h86e333a7_85133007,
        64'h8713fce5_8ce3a1a7,
        64'h8513a007_871367ad,
        64'h06b7f663_08f58c63,
        64'h70070793_67250ab7,
        64'h746304e5_8f637006,
        64'h8713668d_8082852e,
        64'h12f58563_51b00513,
        64'h50000793_00f58963,
        64'h71a00513_70000793,
        64'h0ef58e63_60000793,
        64'h08b7f963_10f58e63,
        64'h30000793_06b76c63,
        64'h80078713_12070963,
        64'h8005871b_04b76263,
        64'h0ee58a63_20078713,
        64'h67858082_01414505,
        64'h18e7a723_47050000,
        64'h27976402_60a2cb3f,
        64'hf0ef1da5_05131d65,
        64'h85930b50_06130000,
        64'h35170000_35978082,
        64'h01414505_1ae7ad23,
        64'h47050000_27976402,
        64'h60a2cdff_f0ef2065,
        64'h05132025_85930b40,
        64'h06130000_35170000,
        64'h3597b791_472df406,
        64'hd5e34705_02579693,
        64'hf406cae3_47350267,
        64'h9693b781_dffff0ef,
        64'h0c800513_f4e796e3,
        64'h8ff54000_0737c000,
        64'h06b7541c_80820141,
        64'h45056402_60a2b709,
        64'h00f60023_47c18082,
        64'h014100e7_90232000,
        64'h07139381_22d71b23,
        64'h17820000_271746cd,
        64'h00071023_27919301,
        64'h00069023_17029281,
        64'h03a7871b_168200c7,
        64'h10233ff6_061b0387,
        64'h869b9301_767d1702,
        64'h00c69023_0367871b,
        64'h92811682_0347869b,
        64'h640260a2_405c00e7,
        64'h80239381_17820287,
        64'h879b4761_405c00e7,
        64'h80239381_17820297,
        64'h879beff0_0613405c,
        64'h0a06d563_02779693,
        64'h473d541c_e9416540,
        64'h10ef8522_a8058593,
        64'h000625b7_0af70663,
        64'h47890364_470300f6,
        64'h80239281_d41047bd,
        64'h16820296_869b4310,
        64'h930102f4_0b230ff7,
        64'hf7931702_0406871b,
        64'h0007d783_93811782,
        64'h0fe6879b_ffed8b85,
        64'h00074783_93011702,
        64'h02f6871b_405400e7,
        64'h80239381_178202f7,
        64'h879b4705_405cf19f,
        64'hf0ef3e80_05130006,
        64'h002310e7_80639201,
        64'h47090ff7_f7930604,
        64'h38230604_22231602,
        64'hd4780296_061b4719,
        64'h0007d783_938102e4,
        64'h00231782_0fe6079b,
        64'h0205c703_cc58cc14,
        64'hc8480104_28230114,
        64'h2623d05c_c0500064,
        64'h10231117_879b1111,
        64'h17b7c41c_4d9449c8,
        64'h0105a803_00c5a883,
        64'h0005d303_4dd8842a,
        64'h459c1c05_8c633807,
        64'ha5230000_27971a05,
        64'h0c63e022_e4061141,
        64'h8082f1a5_05130000,
        64'h25178082_f4850513,
        64'h00002517_808200e7,
        64'h83634501_0247d783,
        64'hf3878793_00002797,
        64'h02a78163_872af467,
        64'hd7830000_27978082,
        64'hfea7ede3_8f99ff86,
        64'hb7830200_c6b702f5,
        64'h05330280_0793fee7,
        64'h8ee3ff86_b7030200,
        64'hc6b7ff87_b7830200,
        64'hc7b78082_ff87b503,
        64'h0200c7b7_80826125,
        64'h70a2a1bf_f0efe43a,
        64'hecc6e8c2_e4bef406,
        64'h72c50513_567d080c,
        64'h86b21838_ec2ee0ba,
        64'hfc36ffff_f517e82a,
        64'h711da43f_f06f72e5,
        64'h0513ffff_f51785aa,
        64'h862e86b2_87368082,
        64'h610560e2_a5dff0ef,
        64'hec06a645_0513002c,
        64'h567d872e_00000517,
        64'h86aa1101_80826161,
        64'h60e2a7bf_f0efe43a,
        64'he4c6e0c2_fc3eec06,
        64'h10387745_0513f83a,
        64'hfffff517_85aa862e,
        64'h86b2f436_715d8082,
        64'h616160e2_aa5ff0ef,
        64'he43ae4c6_e0c2fc3e,
        64'hec067a25_05131018,
        64'h567df83a_f032ffff,
        64'hf51785aa_86aef436,
        64'h715d8082_612560e2,
        64'had1ff0ef_e43aecc6,
        64'he8c2e4be_ec06ae65,
        64'h0513567d_1038858a,
        64'he0baf832_f42e0000,
        64'h051786aa_fc36711d,
        64'hb31d4809_b32d4821,
        64'hbb1d4841_0206e693,
        64'hbb498da2_99020250,
        64'h051385d2_866e86ce,
        64'h001d8413_b7d58622,
        64'h2c859902_00160413,
        64'h02000513_85d286ce,
        64'hbb6d8db2_8aea018c,
        64'he563c019_fc089de3,
        64'hfff8869b_fe0a82e3,
        64'hc51901b7_06330007,
        64'h450378a2_77029902,
        64'h85d286ce_f83af03a,
        64'hf4460705_88b6b7e1,
        64'h78c28df2_8cc27762,
        64'h7e027822_99020200,
        64'h051385d2_86ce866e,
        64'hf072f442_f846fc3a,
        64'h001d8e13_b7c90785,
        64'ha08140ed_8db38cc2,
        64'h018ce863_001c881b,
        64'he4110006_841b8a89,
        64'h00060c9b_8666011c,
        64'hf3638646_000a8863,
        64'h40e78cbb_2a814006,
        64'hfa9302f6_1b63c199,
        64'h0007c583_87ba00f7,
        64'h06339381_02089793,
        64'h00088563_57fd000a,
        64'hb703008a_8d13b7cd,
        64'h8ca22b05_99020200,
        64'h051385d2_86ce001c,
        64'h84138666_b5598de6,
        64'h8aea018b_6563c019,
        64'h9902001d_8c93008a,
        64'h8d1385d2_866e86ce,
        64'h000ac503_ff8764e3,
        64'h001d8d13_00170b1b,
        64'h8dea875a_99020200,
        64'h051385d2_86ce866e,
        64'ha8094705_e00d4b05,
        64'h0006841b_8a89b7ed,
        64'h8f7d67e2_dbe50807,
        64'hf793b769_93014781,
        64'he062e436_17020ff7,
        64'h7713ca09_000aa703,
        64'h0407f613_b755e062,
        64'he4364781_000ab703,
        64'hc7191007_f713bde5,
        64'h4781e062_e436000a,
        64'hb703c719_bff1000a,
        64'ha783b7cd_000a9783,
        64'hc7810807_f793bfd9,
        64'h40e6073b_93fde062,
        64'he43600e7_c63341f7,
        64'hd71b000a_c783cf09,
        64'h0406f713_b789bb7f,
        64'hf0ef854a_85d2866e,
        64'h86ce93fd_40e60733,
        64'h00f74633_43f7d713,
        64'he062e436_000ab783,
        64'hc31d87b6_1006f713,
        64'hb5dd0780_0793eef5,
        64'h09e30750_0793a89d,
        64'h4841e03e_e436008a,
        64'h8413000a_b70347c1,
        64'h0216e693_d4f51ae3,
        64'h07000793_f0f50ce3,
        64'h06f00793_02a7e563,
        64'h12f50f63_07300793,
        64'hb71d0640_07930ef5,
        64'h06630630_0793bddd,
        64'h0c06e693_8082614d,
        64'h6da66d46_6ce67c06,
        64'h7ba67b46_7ae66a0a,
        64'h69aa694a_64ea000d,
        64'h851b740a_70aa9902,
        64'h450185d2_86cefff9,
        64'h8613013d_e463866e,
        64'hda0517e3_0004c503,
        64'h8aa28daa_cf5ff0ef,
        64'h854a85d2_866e86ce,
        64'h93fd40e6_073300f7,
        64'h463343f7_d713e062,
        64'he436000a_b783cf45,
        64'h10c51c63_06400613,
        64'h00c50663_008a8413,
        64'h02085813_270187b6,
        64'h06900613_18022006,
        64'hf7139af9_c3914006,
        64'hf7939acd_00f50363,
        64'h06400793_00f50763,
        64'h48299abd_06900793,
        64'h2ef50463_06200793,
        64'h2ef50663_06f00793,
        64'h2ef50663_05800793,
        64'h2ef50c63_07800793,
        64'he4f514e3_05800793,
        64'h2ef50863_02500793,
        64'h0ca7ef63_00f50c63,
        64'h06200793_0ea7ec63,
        64'h02f50263_00170493,
        64'h06900793_00074503,
        64'h0806e693_0ef60e63,
        64'h0014c603_a0390024,
        64'h87133006_e693a821,
        64'h1006e693_00f60563,
        64'h0014c603_b7e907a0,
        64'h061300c7_89630740,
        64'h0613bf65_84babf75,
        64'h8abe0489_28814881,
        64'h0008d363_008a8793,
        64'h000aa883_00f61d63,
        64'h02a00793_a8998726,
        64'h04c78063_06a00613,
        64'h04c78c63_06800613,
        64'h02f66d63_04c78663,
        64'h00148713_06c00613,
        64'h0004c783_fef671e3,
        64'h0ff7f793_fd07079b,
        64'h00148593_0004c703,
        64'h00e888bb_fd08889b,
        64'h84ae031b_88bbb775,
        64'h84b28aba_40f00c3b,
        64'h0026e693_0007d663,
        64'h00078c1b_008a8713,
        64'h000aa783_fce796e3,
        64'h4c0102a0_0713a825,
        64'h462584ba_06f5ee63,
        64'h4006e693_0ff7f793,
        64'hfd06079b_00148713,
        64'h45a50014_c60306f7,
        64'h17634881_02e00793,
        64'h0004c703_fef671e3,
        64'h0ff7f793_fd07079b,
        64'h00148593_0004c703,
        64'h00e30c3b_fd03031b,
        64'h84ae038b_833bbf75,
        64'h0106e693_b7c90086,
        64'he693b7e1_0046e693,
        64'hb7f90026_e693a025,
        64'h46254c01_06e5e963,
        64'h45a50ff7_7713fd07,
        64'h871b02a7_856302b7,
        64'h8463fcf7_6fe302e7,
        64'h85630014_86130004,
        64'hc78384b2_0016e693,
        64'h02879163_03000413,
        64'h02878f63_02d00413,
        64'ha8210230_05130200,
        64'h059302b0_07134681,
        64'ha15585d2_866e86ce,
        64'h001d8413_00f50863,
        64'h04850250_0793ac81,
        64'h4ba9ec3e_4d81fffb,
        64'h07936b41_cc890913,
        64'h00000917_e589892a,
        64'h8aba84b6_89b28a2e,
        64'he4eee8ea_ece6f0e2,
        64'hf4def8da_f122f506,
        64'hfcd6e152_e54ee94a,
        64'hed267171_808298df,
        64'hf06fc119_b7e1006e,
        64'h033b8082_616160a6,
        64'hd17ff0ef_887e1018,
        64'h0008089b_e43ae876,
        64'he0464746_fc579de3,
        64'hc319fe6f_0fa39f3e,
        64'h0ff37313_02010f13,
        64'h07850307_57330303,
        64'h031b03e3_ee630fff,
        64'h73130307_7f330200,
        64'h0293ff63_0e1b43a5,
        64'h47810410_0313000e,
        64'h04630610_0313020e,
        64'hfe13c721_47810003,
        64'h0463400e_f313fefe,
        64'hfe93e319_4ee68fbe,
        64'he486715d_b7e1006e,
        64'h033b8082_616160a6,
        64'hd97ff0ef_887e1018,
        64'h0008089b_e43ae876,
        64'he0464746_fc579de3,
        64'hc319fe6f_0fa39f3e,
        64'h0ff37313_02010f13,
        64'h07850307_57330303,
        64'h031b03e3_ee630fff,
        64'h73130307_7f330200,
        64'h0293ff63_0e1b43a5,
        64'h47810410_0313000e,
        64'h04630610_0313020e,
        64'hfe13c721_47810003,
        64'h0463400e_f313fefe,
        64'hfe93e319_4ee68fbe,
        64'he486715d_b7a98622,
        64'h9b020016_04130200,
        64'h051385de_86e2b791,
        64'h9b0285de_86e20009,
        64'h4503b7ed_41540cb3,
        64'h02095913_02099913,
        64'hbf89ff27_e3e3009c,
        64'h87b384ea_00148d13,
        64'h67229b02_e43a0200,
        64'h051385de_86e28626,
        64'hb7ad00d6_00230087,
        64'h0633da3d_0087f613,
        64'hbf9d02b0_06130087,
        64'h06b3c611_0047f613,
        64'hbfa10620_06130087,
        64'h06b3f886_ece346fd,
        64'hf6d898e3_4689b7bd,
        64'h05800613_008706b3,
        64'hfa86e7e3_46fd8082,
        64'h61658532_6d426ce2,
        64'h7c027ba2_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_0b37e163,
        64'h415607b3_0209d993,
        64'h1982000a_09630094,
        64'h06330b2c_9663197d,
        64'h412d0633_01248d33,
        64'hfff70c93_00870933,
        64'hcbcd84d6_8b8d0405,
        64'h00c68023_02d00613,
        64'h008706b3_08080463,
        64'h00d40b63_02000693,
        64'h040500c6_80230300,
        64'h06130087_06b30286,
        64'he66346fd_040500c6,
        64'h80230780_06130087,
        64'h06b30486_e06346fd,
        64'head10207_f6930ad8,
        64'h966346c1_4401bf55,
        64'hfe6e0fa3_00870e33,
        64'h0405a0e9_02c89a63,
        64'h84364609_02c88163,
        64'h14794641_c285fff4,
        64'h06930286_95639281,
        64'h02099693_00868763,
        64'h92811682_cc0dee15,
        64'h4007f613_ca3d0107,
        64'hf61302b4_1e6300a4,
        64'h7463c609_03000313,
        64'h02000593_91010209,
        64'h9513fea4_69e3fe6e,
        64'h0fa30087_0e330405,
        64'h00b40963_a8010300,
        64'h03130200_05939101,
        64'h02069513_39fdc191,
        64'h00c7f593_00081563,
        64'hc6190009_89630017,
        64'hf613040a_1a6359e6,
        64'h56c68ab2_8bae8b2a,
        64'h8c362a01_e86aec66,
        64'he8caeca6_f486f062,
        64'hf45ef85a_fc560027,
        64'hfa13e4ce_e0d2478a,
        64'h843ef0a2_71598082,
        64'h8302658c_0005b303,
        64'hc5098082_808200a5,
        64'h802395b2_00d67563,
        64'hbbe102f0_00efd3e5,
        64'h05130000_4517bd35,
        64'hb0250513_85a60000,
        64'h45170470_00efaf65,
        64'h05130000_4517cd09,
        64'h84aada9f_f0ef8552,
        64'h865a020a_a5830630,
        64'h00efd5a5_05130000,
        64'h4517f579_90e30804,
        64'h84930770_00ef2985,
        64'ha4850513_00004517,
        64'hff2c17e3_089000ef,
        64'h0905cfa5_05130000,
        64'h45170009_45830704,
        64'h8c130284_89130a30,
        64'h00efd825_05130000,
        64'h45170af0_00efd765,
        64'h05130000_4517708c,
        64'h0bd000ef_d6c50513,
        64'h00004517_6c8c0cb0,
        64'h00efd625_05130000,
        64'h4517688c_ff2c17e3,
        64'h0dd000ef_0905d4e5,
        64'h05130000_45170009,
        64'h45830109_0c130f30,
        64'h00efd6a5_05130000,
        64'h4517fe99_17e31030,
        64'h00ef0905_d7450513,
        64'h00004517_00094583,
        64'hff048913_119000ef,
        64'hd6850513_00004517,
        64'h125000ef_d5e50513,
        64'h85ce0000_4517bf15,
        64'hd4a50513_85ce0000,
        64'h451713f0_00efbee5,
        64'h05130000_4517cd09,
        64'h4b910804_89aa8a8a,
        64'hea7ff0ef_850a4605,
        64'h710144ac_161000ef,
        64'hd5850513_00004517,
        64'h45d616f0_00efd465,
        64'h05130000_451745c6,
        64'h17d000ef_d2c50513,
        64'h00004517_65a618b0,
        64'h00efd225_05130000,
        64'h45177582_199000ef,
        64'hd1850513_00004517,
        64'h65e21a70_00efd0e5,
        64'h05130000_451745d2,
        64'h1b5000ef_d0450513,
        64'h00004517_45c21c30,
        64'h00efcfa5_05130000,
        64'h451745b2_1d1000ef,
        64'hcf050513_00004517,
        64'h45a21df0_00efce65,
        64'h05130000_45176582,
        64'h1ed000ef_cd450513,
        64'h00004517_b75554f9,
        64'h1fd000ef_cc450513,
        64'h00004517_fa843583,
        64'h20d000ef_cbc50513,
        64'h00004517_faa43423,
        64'hc11df71f_f0ef848a,
        64'h850a4585_46057101,
        64'h22d000ef_cc450513,
        64'h00004517_80826125,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h64468526_60e6fa04,
        64'h011354fd_259000ef,
        64'hcc850513_00004517,
        64'hc51df39f_f0ef8b2e,
        64'h8a2a1080_e862ec5e,
        64'hf456fc4e_e0cae4a6,
        64'hec86f05a_f852e8a2,
        64'h711d8082_014160a2,
        64'h557d28f0_00efcde5,
        64'h05130000_451785aa,
        64'hc9095600_10efe406,
        64'hc0c50513_46051141,
        64'h00003517_86aab76d,
        64'h45012b70_00efce65,
        64'h05130000_4517bf6d,
        64'h55752c70_00efcc65,
        64'h05130000_4517c909,
        64'h85aa1500_10ef8522,
        64'hbfd15579_2e1000ef,
        64'hcb850513_00004517,
        64'hc90985aa_441000ef,
        64'h852285aa_c5c40413,
        64'h00003417_41508082,
        64'h01416402_60a2557d,
        64'h30d000ef_cc450513,
        64'h00004517_ed014350,
        64'h00ef4501_321000ef,
        64'he022e406_cc650513,
        64'h11410000_45178082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_00a78223,
        64'h0ff57513_00d78023,
        64'h0085551b_0ff57693,
        64'h00d78623_f8000693,
        64'h00078223_01e71793,
        64'h470d02b5_553b0045,
        64'h959b8082_00a78023,
        64'hdf650207_77130147,
        64'hc70307fa_478d8082,
        64'h02057513_0147c503,
        64'h07fa478d_80820005,
        64'h45038082_00b50023,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_100004b7,
        64'h18858593_00003597,
        64'hf1402573_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_3e7020ef,
        64'h40000137_03249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
