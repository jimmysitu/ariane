/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 2095;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00000078_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000078_36313025,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000078_36313025,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_78323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000a64_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h00000a64_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_0000000a,
        64'h78363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h0000000a_78363130,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h0000000a_78363130,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_00000a64,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_00000a64,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_00000a64,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_00000a64,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h00000000_00000a78,
        64'h25202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h0000000a_21206465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_0a212064,
        64'h656c6961_66206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a2120,
        64'h64656c69_61662067,
        64'h69666e6f_43204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_002e2e2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd0080000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h08090000_38000000,
        64'hda0b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_a001830f,
        64'he0ef1e25_05130000,
        64'h15178402_5dc58593,
        64'h00000597_10000437,
        64'he901dcaf_d0ef1000,
        64'h053765a1_856fe0ef,
        64'h20050513_00001517,
        64'h950fe0ef_24040513,
        64'h86afe0ef_21450513,
        64'h00001517_964fe0ef,
        64'h24040513_000f4437,
        64'h882fe0ef_20450513,
        64'h00001517_d56fd0ef,
        64'he022e406_a0050513,
        64'h20058593_11410262,
        64'h653765f1_80820141,
        64'h421c9201_00f69023,
        64'h16024789_26416402,
        64'h60a28082_01414505,
        64'h640260a2_80820141,
        64'h450500f6_10233ff7,
        64'h879b9201_77fd1602,
        64'h640260a2_0326061b,
        64'hfe0756e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d783ef9d,
        64'ha0119281_16820306,
        64'h069b4050_e129de0f,
        64'he0ef842a_e406e022,
        64'h60000593_4681862e,
        64'h11418082_0141439c,
        64'h938100e6_90231782,
        64'h47090106_079b6402,
        64'h60a28082_01414505,
        64'h64e7af23_47050000,
        64'h07976402_60a2948f,
        64'he0ef64a5_051365e5,
        64'h859335c0_06130000,
        64'h15170000_15978082,
        64'h01414505_640260a2,
        64'h80820141_450568e7,
        64'haa234705_00000797,
        64'h640260a2_97efe0ef,
        64'h68050513_69458593,
        64'h35d00613_00001517,
        64'h00001597_80820141,
        64'h450500e7_90233ff7,
        64'h071b9381_777d1782,
        64'h640260a2_0326079b,
        64'hfe0756e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d783ebd9,
        64'ha0119281_16820306,
        64'h069b4050_e53deb0f,
        64'he0ef70e7_97238522,
        64'h80058593_46014685,
        64'h47450000_07976585,
        64'hc0dfe0ef_85224585,
        64'h00e79023_93811782,
        64'h2791862e_20000713,
        64'h405cfee7_9de30785,
        64'h00078023_08d61263,
        64'h20058713_87ae842a,
        64'h11168693_7407a623,
        64'h111116b7_00000797,
        64'h5150c979_e022e406,
        64'h11418082_0141853e,
        64'h478576e7_a4234705,
        64'h00000797_640260a2,
        64'ha52fe0ef_75450513,
        64'h76858593_32c00613,
        64'h00001517_00001597,
        64'h80820141_853e00a0,
        64'h37b36402_60a2f50f,
        64'he0efa005_85934601,
        64'h46818522_65adf17d,
        64'h4785f64f_e0ef7005,
        64'h85934681_658d4930,
        64'h80820141_853e6402,
        64'h60a24785_7ce7a523,
        64'h47050000_0797ab0f,
        64'he0ef7b25_05137c65,
        64'h859332d0_06130000,
        64'h15170000_159702f7,
        64'h0963842a_11178793,
        64'h111117b7_7e07ad23,
        64'h51580000_0797cd25,
        64'he022e406_1141bd85,
        64'hbd8fe0ef_4505dc07,
        64'h80e30807_f7930007,
        64'hd783b3f1_450582e7,
        64'ha2234705_00001797,
        64'hb0afe0ef_80c50513,
        64'h82058593_48e00613,
        64'h00002517_00002597,
        64'hb7e9ffcf_e0ef85d2,
        64'hfd3798e3_852285ca,
        64'h46014685_03444783,
        64'hc0a1c329_04077713,
        64'h0007d703_93811782,
        64'h03e7879b_405ce205,
        64'h10e30ff4_f49334fd,
        64'h833fe0ef_a01d300a,
        64'h0a134985_c54fe0ef,
        64'h00e79023_04076713,
        64'h02800493_500a0913,
        64'h0007d703_93818ad7,
        64'h142346c1_00001717,
        64'h178200d7_102303e7,
        64'h879b9301_17020047,
        64'h871b4505_6a05405c,
        64'h04000693_00f70463,
        64'h08000693_478d0374,
        64'h470308f7_1b631117,
        64'h87931111_17b78e07,
        64'ha2235058_00001797,
        64'hbd694505_d939c63f,
        64'hf0ef8522_50058593,
        64'hdc1c0319_75b75007,
        64'h879b0319_77b700f6,
        64'h90234789_bd7d4505,
        64'hdd2dc87f_f0ef8522,
        64'h08058593_dc1c02fa,
        64'hf5b70807_879b02fa,
        64'hf7b700f6_90234789,
        64'hb5a5fe07_56e38b89,
        64'h4107571b_0107971b,
        64'h93c117c2_0006d783,
        64'hef9da011_92811682,
        64'h0306069b_4050f005,
        64'h14e3915f_e0ef6000,
        64'h05931006_06134681,
        64'h03b90637_b5f5439c,
        64'h93811782_27c1405c,
        64'h00e78023_00476713,
        64'h0007c703_93811782,
        64'h0287879b_4501405c,
        64'hd60fe0ef_3e800513,
        64'h0af70a63_479d5478,
        64'hf921d17f_f0ef8522,
        64'h00f69023_47895c0c,
        64'hb5e5fe07_56e38b89,
        64'h4107571b_0107971b,
        64'h93c117c2_0006d783,
        64'hefc9a011_92811682,
        64'h0306069b_4050f159,
        64'h993fe0ef_9ee79823,
        64'h85226000_05931645,
        64'h46854745_00001797,
        64'h81000637_ef1fe0ef,
        64'h458500e7_90239381,
        64'h17822791_860a0400,
        64'h0713415c_80826165,
        64'h45056a06_69a66946,
        64'h64e6a2e7_a0234705,
        64'h00001797_740670a6,
        64'hd0afe0ef_a0c50513,
        64'ha2058593_1f300613,
        64'h00002517_00002597,
        64'h80826165_6a0669a6,
        64'h694664e6_740670a6,
        64'h4505d135_a0ffe0ef,
        64'h85226000_05934681,
        64'h20060613_dd1c03b9,
        64'h06372007_879b0beb,
        64'hc7b78082_61656a06,
        64'h69a66946_64e67406,
        64'h70a64505_a8e7a523,
        64'h47050000_1797d70f,
        64'he0efa725_0513a865,
        64'h85931f40_06130000,
        64'h25170000_25978082,
        64'h61654505_6a0669a6,
        64'h694664e6_00f61023,
        64'h3ff7879b_920177fd,
        64'h16027406_70a60326,
        64'h061bfe07_55e38b89,
        64'h4107571b_0107971b,
        64'h93c117c2_0006d783,
        64'h12079a63_a0199281,
        64'h16820306_069b4050,
        64'he145aadf_e0ef8522,
        64'h60000593_46811006,
        64'h0613dd1c_03b90637,
        64'h5007879b_031977b7,
        64'h0af70163_479d5578,
        64'h1ae78863_470910e7,
        64'h8b634705_03454783,
        64'h08f71363_842a1117,
        64'h87931111_17b7b207,
        64'hae235158_00001797,
        64'h10050263_fc02f802,
        64'hf402f002_ec02e802,
        64'he402e002_e0d2e4ce,
        64'he8caeca6_f0a2f486,
        64'h71598082_01414505,
        64'hb6e7a723_47050000,
        64'h179760a2_e56fe0ef,
        64'hb5850513_b6c58593,
        64'h2b700613_00002517,
        64'h00002597_b75d00c6,
        64'h90239241_16428e5d,
        64'h06228fd9_0017e793,
        64'h820503f7_f793071a,
        64'h00965713_0006d783,
        64'hfee5e8e3_27859241,
        64'h03079613_02f8573b,
        64'hf8a78be3_a0197ff0,
        64'h05134785_80820141,
        64'h00f69023_0047e793,
        64'h450160a2_0006d783,
        64'hdfed8b89_0006d783,
        64'h00e69023_93411742,
        64'h8f5d0017_e7930ff7,
        64'hf7930722_83050006,
        64'hd783bfd9_c0e7a523,
        64'h47050000_1797ef0f,
        64'he0efbf25_0513c065,
        64'h85932b80_06130000,
        64'h25170000_25978082,
        64'h01414505_60a2f675,
        64'h93410305_171302f5,
        64'hfc63367d_0017151b,
        64'h02e857bb_07178e63,
        64'h03654783_00f69023,
        64'h93c117c2_9be993c1,
        64'h17c24705_46250006,
        64'hd7839281_168202c6,
        64'h869b4889_00852803,
        64'h415404f7_18631117,
        64'h87931111_17b7c807,
        64'ha2235158_00001797,
        64'h10050063_e4061141,
        64'h80820141_439c9381,
        64'h00e69023_17824709,
        64'h0106079b_640260a2,
        64'h80820141_4505cae7,
        64'haa234705_00001797,
        64'h640260a2_f9efe0ef,
        64'hca050513_cb458593,
        64'h19f00613_00002517,
        64'h00002597_80820141,
        64'h45056402_60a28082,
        64'h01414505_cee7a523,
        64'h47050000_17976402,
        64'h60a2fd4f_e0efcd65,
        64'h0513cea5_85931a00,
        64'h06130000_25170000,
        64'h25978082_01414505,
        64'h00e79023_3ff7071b,
        64'h9381777d_17826402,
        64'h60a20326_079bfe07,
        64'h56e38b89_4107571b,
        64'h0107971b_93c117c2,
        64'h0006d783_ebd9a011,
        64'h92811682_0306069b,
        64'h4050e53d_d07fe0ef,
        64'hd6e79223_85226000,
        64'h05931641_46854745,
        64'h00001797_01000637,
        64'ha64ff0ef_85224585,
        64'h00e79023_93811782,
        64'h2791862e_04000713,
        64'h405cfee7_9de30785,
        64'h00078023_08d61363,
        64'h04058713_87ae842a,
        64'h11168693_da07a223,
        64'h111116b7_00001797,
        64'h5150cd61_e022e406,
        64'h1141b765_00e69023,
        64'h00476713_9b619341,
        64'h17420006_d7039281,
        64'h168203e7_869b405c,
        64'hb5fd4505_d551d91f,
        64'he0ef8522_60058593,
        64'h46094681_02f40ba3,
        64'h65a14789_f00515e3,
        64'hdabfe0ef_85227005,
        64'h85934681_658d4830,
        64'hb7a94501_439c9381,
        64'h178227c1_405c04f7,
        64'h01634791_547800e7,
        64'h80230ff7_77130206,
        64'he71300c5_94630026,
        64'he7130ff6_f6930007,
        64'hc6839381_17820287,
        64'h879b460d_03744583,
        64'h405ca13f_e0ef3e80,
        64'h051300f6_90234789,
        64'hb7256007_8613f2e6,
        64'h98e32007_86134711,
        64'h02e40ba3_03b707b7,
        64'h470df2f7_18e347a1,
        64'h48588082_01414505,
        64'he6e7af23_47050000,
        64'h17976402_60a2969f,
        64'he0efe6a5_0513e7e5,
        64'h85931120_06130000,
        64'h25170000_2597b7e5,
        64'hf4e7e1e3_4501478d,
        64'h4958b749_50078613,
        64'h80820141_640260a2,
        64'h4505ece7_a0234705,
        64'h00001797_9a7fe0ef,
        64'hea850513_ebc58593,
        64'h11300613_00002517,
        64'h00002597_80820141,
        64'h640260a2_450500f6,
        64'h10233ff7_879b9201,
        64'h77fd1602_0326061b,
        64'hfe0756e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d783e3e1,
        64'ha0119281_16820306,
        64'h069b4050_ed05ed9f,
        64'he0ef8522_60000593,
        64'h468106e6_8f631007,
        64'h86134711_02e40ba3,
        64'h03b707b7_47090ce7,
        64'h88635474_07522000,
        64'h57378ff9_17820ff7,
        64'h879300ff_07b77818,
        64'h14f70e63_47850344,
        64'h47030af7_0e634789,
        64'h03654703_08f71a63,
        64'h842a1117_87931111,
        64'h17b7f807_a0235158,
        64'h00001797_c565e022,
        64'he4061141_b7a9439c,
        64'h938100e6_90231782,
        64'h47090106_079b8082,
        64'h61054505_64a2fae7,
        64'ha6234705_00001797,
        64'h644260e2_a97fe0ef,
        64'hf9850513_fac58593,
        64'h0b900613_00002517,
        64'h00002597_bfb14505,
        64'h00e79023_3ff7071b,
        64'h9381777d_17820326,
        64'h079bfe07_56e38b89,
        64'h4107571b_0107971b,
        64'h93c117c2_0006d783,
        64'hefb1a011_92811682,
        64'h0306069b_4050f951,
        64'hfc3fe0ef_02e79023,
        64'h85223005_85934601,
        64'h46854745_00001797,
        64'h65add1ef_f0ef8522,
        64'h458500e7_90239381,
        64'h17822791_86264721,
        64'h405c8082_610564a2,
        64'h644260e2_450504e7,
        64'ha6234705_00001797,
        64'hb33fe0ef_03450513,
        64'h04858593_0ba00613,
        64'h00002517_00002597,
        64'h80826105_64a26442,
        64'h60e24505_cd15830f,
        64'hf0ef8522_70058593,
        64'h4681658d_4830fee7,
        64'h9de30785_00078023,
        64'h02d61663_00858713,
        64'h87ae84ae_842a1116,
        64'h86930a07_a5231111,
        64'h16b70000_17975150,
        64'hc17de426_e822ec06,
        64'h11018082_61054505,
        64'h64a20ce7_a4234705,
        64'h00001797_644260e2,
        64'hbb3fe0ef_0b450513,
        64'h0c858593_07e00613,
        64'h00002517_00002597,
        64'hb7650097_90234318,
        64'h93818cf5_93011782,
        64'h17022791_0107871b,
        64'h16fd6685_405cf171,
        64'h8c2ff0ef_65854681,
        64'h862e84ae_bfc910e7,
        64'hae234705_00001797,
        64'hc03fe0ef_10450513,
        64'h11858593_07f00613,
        64'h00002517_00002597,
        64'h80826105_64a26442,
        64'h60e24505_cb8d3037,
        64'hf793439c_93811782,
        64'h0247879b_415c02f7,
        64'h1163842a_11178793,
        64'h111117b7_1607a523,
        64'h51580000_1797c541,
        64'he426e822_ec061101,
        64'hb6c14905_ea0501e3,
        64'h1f8000ef_8522b6f9,
        64'h4905eaf7_08e34789,
        64'h0b94c703_b5c1c407,
        64'h9de30a24_c78300e7,
        64'h8e634711_bcd713e3,
        64'h0b94c703_bd3902f4,
        64'h0e234785_d85fe0ef,
        64'h00e79023_00476713,
        64'h3e800513_0007d703,
        64'hb9014905_def709e3,
        64'h47850b94_c703be05,
        64'h1ce32850_00ef8522,
        64'h85a6c005_12e36880,
        64'h00ef8522_d47c4795,
        64'hbfd59341_17420007,
        64'hd703eb15_8b099341,
        64'h17420007_d70300e7,
        64'h90230017_67130007,
        64'hd7039381_178202c7,
        64'h879bc207_0ee38b21,
        64'h00075703_93011702,
        64'h03e7871b_405cdfff,
        64'he0ef00e7_90230087,
        64'h67130007_d70300e6,
        64'h90239381_93411742,
        64'h9b699341_17421782,
        64'h03e7879b_0006d703,
        64'h92811682_02c7869b,
        64'h38850513_6505405c,
        64'hec079ee3_03c44783,
        64'heef712e3_47a14858,
        64'heee7f6e3_478d00d1,
        64'h4703bfbd_d47c4795,
        64'hfee7f5e3_47850374,
        64'h4703dbed_8b89bba1,
        64'hd3f10a24_c783d47c,
        64'h4799c719_00c7f713,
        64'hb755d47c_479100f9,
        64'hf8630374_4783c30d,
        64'h00c7f713_b311892a,
        64'hb3214905_ee0505e3,
        64'h493000ef_85221005,
        64'h859303a2_05b7ee07,
        64'h9ee30a24_c78312e6,
        64'hfb634685_ffc7871b,
        64'h14e78c63_471d547c,
        64'hd00519e3_39f000ef,
        64'h852285a6_d0051fe3,
        64'h7a2000ef_8522d47c,
        64'h479d06e9_f3630374,
        64'h4703cf21_0307f713,
        64'h0c44c783_d07c8fd9,
        64'h0d44c703_d07c8fd9,
        64'h0087171b_0d54c703,
        64'hd07c2781_8fd90107,
        64'h979b0d64_c783d078,
        64'h0187971b_0d74c783,
        64'hd60515e3_3f7000ef,
        64'h15648493_85221564,
        64'h85930000_1497d805,
        64'h10e33da0_00ef8522,
        64'hbb454905_d9410110,
        64'h00ef8522_d47c4795,
        64'hf8e7ffe3_47850374,
        64'h4703d3dd_8b8900d1,
        64'h4783d7dd_0004c783,
        64'h1007c963_00248783,
        64'hed695ec0_00ef8522,
        64'h858adc05_12e341e0,
        64'h00ef8522_c7918b91,
        64'h0014c783_dc051be3,
        64'h302000ef_852285a6,
        64'hde0511e3_3c3000ef,
        64'h8522bd09_e8f708e3,
        64'h47850344_4703e8f7,
        64'h1de34791_54781efa,
        64'h69630374_4783c789,
        64'h8b890c44_c783d07c,
        64'h8fd90d44_c703d07c,
        64'h8fd90087_171b0d54,
        64'hc703d07c_27818fd9,
        64'h0107979b_0d64c783,
        64'hd0780187_971b0d74,
        64'hc783e205_1ee34c90,
        64'h00ef2284_84938522,
        64'h22848593_00001497,
        64'he40519e3_4ac000ef,
        64'h8522ef3a_1be30364,
        64'h4a03eee7_ffe3478d,
        64'h03544703_bdd9ac05,
        64'h8593dc1c_0121f5b7,
        64'hac07879b_0121f7b7,
        64'hbf8502f4_0a234789,
        64'hbdcd8405_8593dc1c,
        64'h017d85b7_8407879b,
        64'h017d87b7_02f70063,
        64'h47890364_4703ea05,
        64'h14e3de6f_f0ef8522,
        64'hf0d711e3_bdf14905,
        64'hf0f705e3_479500f6,
        64'hf7630ff7_f793fff7,
        64'h079b4685_03444703,
        64'hffed8b89_00074783,
        64'h93011702_02f7071b,
        64'h405800e7_80234709,
        64'h938100d7_10231782,
        64'h3ff6869b_930176fd,
        64'h02f7879b_170200c6,
        64'h90230327_871b9281,
        64'h16820307_869b567d,
        64'h405c02f4_0a234785,
        64'hc949cb4f_f0ef8522,
        64'h10000593_40ff8637,
        64'h4681bf89_490550e7,
        64'haa234705_00001797,
        64'hffbfe0ef_4fc50513,
        64'h4f858593_23f00613,
        64'h00002517_00002597,
        64'hbfa500a0_39333c20,
        64'h00ef8522_20000593,
        64'hf8f705e3_47915478,
        64'h1ee78263_471510e7,
        64'h83634709_19378763,
        64'h49850344_4783fd3d,
        64'h892ad1cf_f0ef8522,
        64'h70000593_46814830,
        64'hf9410e70_00ef8522,
        64'ha8058593_dc1c018c,
        64'hc5b7a807_879b018c,
        64'hc7b7f54d_d55ff0ef,
        64'h852202f5_0a234795,
        64'hfae791e3_8ff54000,
        64'h0737c000_06b7551c,
        64'h8082610d_7a4679e6,
        64'h690a64aa_854a644a,
        64'h60ea4905_5ce7a123,
        64'h47050000_17978a8f,
        64'hf0ef5aa5_05135a65,
        64'h85932400_06130000,
        64'h25170000_2597a01d,
        64'h4905cd69_d9eff0ef,
        64'h85224581_46014681,
        64'h9c0ff0ef_71050513,
        64'h650904f7_0b634789,
        64'h02050e23_dd1ca807,
        64'h879b0006_27b70365,
        64'h470302f5_0a2302f5,
        64'h0ba34785_04f71163,
        64'h842a1117_87931111,
        64'h17b76207_a8235158,
        64'h00001797_10050463,
        64'hfc02f802_f402f002,
        64'hec02e802_e402e002,
        64'h0004b023_9881f8d2,
        64'hfccee14a_e922ed06,
        64'h05f10493_e5267135,
        64'hb5f1d07c_02e40aa3,
        64'h0097d79b_00f6f713,
        64'h0126569b_00e797bb,
        64'h00f6f713_00e797bb,
        64'h27850086_d69b2709,
        64'h8b1d8fcd_42100077,
        64'h571b8fe5_92010167,
        64'h559b1602_00a6979b,
        64'h26812701_01c7861b,
        64'h42944318_42109281,
        64'h93019201_16821702,
        64'h16020187_869b0147,
        64'h871b0107_861bc004,
        64'h8493405c_f00515e3,
        64'he8aff0ef_85229004,
        64'h85934681_64854830,
        64'hfd11e9cf_f0ef3000,
        64'h05931234_0637c83c,
        64'hc4381234_07b7c47c,
        64'hc070c02c_0007d783,
        64'h00075703_00065603,
        64'h0005d583_93819301,
        64'h92019181_17821702,
        64'h16021582_27f10187,
        64'h871b0147_861b0107,
        64'h859b8522_4681405c,
        64'hf535eecf_f0ef8522,
        64'h20000593_46014681,
        64'hd81c4785_00075463,
        64'h02179713_80826105,
        64'h450564a2_74e7ad23,
        64'h47050000_17976442,
        64'h60e2a44f_f0ef7465,
        64'h05137425_85936700,
        64'h06130000_25170000,
        64'h2597b751_f6e798e3,
        64'h8ff54000_0737c000,
        64'h06b7551c_80826105,
        64'h64a26442_60e24505,
        64'h78e7af23_47050000,
        64'h1797a84f_f0ef7865,
        64'h05137825_85936710,
        64'h06130000_25170000,
        64'h25978082_61054505,
        64'h64a26442_60e2d165,
        64'hf82ff0ef_85221000,
        64'h059340ff_86374681,
        64'h0807c863_2781439c,
        64'h93811782_27c1405c,
        64'ha015c911_fa6ff0ef,
        64'h85224581_46014681,
        64'h02075b63_02f79713,
        64'h439c9381_17820247,
        64'h879b405c_cb99445c,
        64'h08f70463_47890365,
        64'h470306f7_1263842a,
        64'h11178793_111117b7,
        64'h8207a723_51580000,
        64'h2797cd4d_e426e822,
        64'hec061101_80826145,
        64'h450169a2_694264e2,
        64'h00f69023_47897402,
        64'h70a2b775_dd25811f,
        64'hf0ef86e7_97238522,
        64'h80058593_864e4685,
        64'h470d0000_27976589,
        64'hb799f4c7_13e30107,
        64'h77334000_0637c000,
        64'h08375518_bff9f406,
        64'h4fe302f7_16134318,
        64'h93011702_0247871b,
        64'h80826145_450569a2,
        64'h694264e2_740270a2,
        64'h00f61023_3ff7879b,
        64'h920177fd_16020326,
        64'h061bfe07_56e38b89,
        64'h4107571b_0107971b,
        64'h93c117c2_0006d783,
        64'he3c1a011_92811682,
        64'h0306069b_4050ed05,
        64'h89bff0ef_8ee79d23,
        64'h85229005_8593864e,
        64'h86a60270_07130000,
        64'h27976589_08f48863,
        64'h4785dfff_f0ef8522,
        64'h85a6864a_e13d79a0,
        64'h00ef2000_059300f7,
        64'h0763842a_89ae8936,
        64'h20000713_439c9381,
        64'h17822791_eb594558,
        64'h0ae80863_415c84b2,
        64'h47090365_4803e44e,
        64'he84af022_f406ec26,
        64'h71798082_61454501,
        64'h421c69a2_694264e2,
        64'h920100f6_90231602,
        64'h47892641_740270a2,
        64'hb775dd25_927ff0ef,
        64'h98e79223_85221005,
        64'h8593864e_4685474d,
        64'h00002797_6585b799,
        64'hf4c713e3_01077733,
        64'h40000637_c0000837,
        64'h5518bff9_f4064fe3,
        64'h02f71613_43189301,
        64'h17020247_871b8082,
        64'h61454505_69a26942,
        64'h64e27402_70a200f6,
        64'h10233ff7_879b9201,
        64'h77fd1602_0326061b,
        64'hfe0756e3_8b894107,
        64'h571b0107_971b93c1,
        64'h17c20006_d783e3c1,
        64'ha0119281_16820306,
        64'h069b4050_ed059b1f,
        64'hf0efa0e7_98238522,
        64'h20058593_864e86a6,
        64'h03700713_00002797,
        64'h658508f4_88634785,
        64'hf15ff0ef_852285a6,
        64'h864ae13d_0b1000ef,
        64'h20000593_00f70763,
        64'h842a89ae_89362000,
        64'h0713439c_93811782,
        64'h2791eb59_45580ae8,
        64'h0863415c_84b24709,
        64'h03654803_e44ee84a,
        64'hf022f406_ec267179,
        64'h808200a8_a02308b7,
        64'h91230208_d8930805,
        64'h051b08e7_902308c7,
        64'ha2231882_02300713,
        64'h97aa0588_889b83f5,
        64'h02069793_026585bb,
        64'h9e3901e7_073b7741,
        64'hff0718e3_07a100ee,
        64'h073b0007_912301d7,
        64'h9023c3d8_6e410210,
        64'h0e938732_01e8083b,
        64'h08050793_00c8083b,
        64'h01071f1b_7841ce85,
        64'hfff7069b_0016871b,
        64'hc3990006_871b93c1,
        64'h17c20107_d69b04e8,
        64'h69630007_881b4681,
        64'h02b307bb_00f37333,
        64'h26016741_0007d783,
        64'h93811782_0048879b,
        64'h137d6305_00452883,
        64'h80820141_00a03533,
        64'h60a2acdf_f0efe406,
        64'h70000593_46811141,
        64'h4930b339_d07c0097,
        64'hd79b00f7_17bb00f6,
        64'h779300f7_173b0086,
        64'h561b2705_27898b9d,
        64'h8f550077_d79b8f65,
        64'h0167d69b_c0048493,
        64'h00a6171b_b381d07c,
        64'h00a7979b_278593a9,
        64'h178ad4d7_18e34685,
        64'hcb198b0d_0166d71b,
        64'h26010007_079b4394,
        64'h42904318_93019381,
        64'h92814210_17821682,
        64'h17029201_27f11602,
        64'h0187869b_0147871b,
        64'h0107861b_405cd405,
        64'h1be3b5df_f0ef8522,
        64'h90048593_46816485,
        64'hb59902f4_0aa34789,
        64'hbb854505_d16db79f,
        64'hf0ef8522_30000593,
        64'h46014681_ee19c830,
        64'h8e654390_93811782,
        64'h27c1405c_a809c47c,
        64'hc438c074_c0300007,
        64'hd7830007_57030006,
        64'hd6830006_56039381,
        64'h93019281_92011782,
        64'h17021682_160227f1,
        64'h0187871b_0147869b,
        64'h0107861b_74c1405c,
        64'hdc0518e3_bd7ff0ef,
        64'h85222000_05934601,
        64'h4681de04_91e3fed7,
        64'h9ee38ff1_431c00d7,
        64'h86638ff1_431c9301,
        64'h17020247_071b01f0,
        64'h06b701f0_06374058,
        64'h821ff0ef_00f71023,
        64'h0047e793_3e800513,
        64'h00075783_dfed8b89,
        64'h00075783_00f71023,
        64'h0017e793_00075783,
        64'h93010207_971302c7,
        64'h879be207_0de38b21,
        64'h00075703_93011702,
        64'h03e7871b_405c867f,
        64'hf0ef00f6_90230087,
        64'he7933885_05136505,
        64'h0006d783_928100f7,
        64'h102393c1_17c29be9,
        64'h93c117c2_168203e6,
        64'h869b0007_57839301,
        64'h170202c6_871bfff5,
        64'h8ff1431c_c7818ff1,
        64'h431c9301_17020246,
        64'h871b84aa_01f00637,
        64'h4054ca5f_f0ef8522,
        64'hb0058593_46014681,
        64'h02f40e23_65854785,
        64'h0c075d63_02779713,
        64'hd8184705_00075463,
        64'h02179713_bf7541ff,
        64'h8637fd47_92e3485c,
        64'hfd3795e3_40ff8637,
        64'h85220364_4783ee05,
        64'h13e385a6_4681cf1f,
        64'hf0ef8522_460185ca,
        64'h46810207_c9632781,
        64'h439c9381_178227c1,
        64'h405cf005_15e3d11f,
        64'hf0efa829_90048493,
        64'h4a214989_70090913,
        64'h64ad690d_02f40aa3,
        64'h47851af7_0f631aa0,
        64'h0713431c_93011702,
        64'h27414058_80826145,
        64'h45056a02_69a26942,
        64'h64e2d8e7_ac234705,
        64'h00002797_740270a2,
        64'h883ff0ef_d8450513,
        64'hd8058593_16100613,
        64'h00003517_00003597,
        64'hb785f4e7_96e38ff5,
        64'h40000737_c00006b7,
        64'h551ca0a9_ffed8b89,
        64'h0006c783_92811682,
        64'h02f7069b_405800a7,
        64'h80239381_178202f7,
        64'h879b405c_faf512e3,
        64'h4789c925_dafff0ef,
        64'h85228005_85931aa0,
        64'h06134681_65858082,
        64'h61456a02_69a26942,
        64'h64e27402_70a24505,
        64'he0e7af23_47050000,
        64'h2797905f_f0efe065,
        64'h0513e025_85931620,
        64'h06130000_35170000,
        64'h35978082_61456a02,
        64'h69a26942_64e27402,
        64'h70a24505_c521e09f,
        64'hf0ef8522_45814601,
        64'h46810007_596302f7,
        64'h9713439c_93811782,
        64'h0247879b_405ccb99,
        64'h445c0af7_06634789,
        64'hc95c4791_03654703,
        64'h04f71563_842a1117,
        64'h87931111_17b7e807,
        64'haa235158_00002797,
        64'hc16de052_e44ee84a,
        64'hec26f022_f4067179,
        64'hb76900e7_90232501,
        64'h3ff7071b_777d4509,
        64'he311ffe5_77139141,
        64'h15420007_d5039381,
        64'h02051793_0325051b,
        64'h80826105_45056902,
        64'h64a2eee7_a0234705,
        64'h00002797_644260e2,
        64'h9cbff0ef_ecc50513,
        64'hec858593_44b00613,
        64'h00003517_00003597,
        64'hb76d00f6_10230200,
        64'h0793d6dd_0206f693,
        64'h00065683_80826105,
        64'h690264a2_644260e2,
        64'h4505f2e7_a4234705,
        64'h00002797_a0fff0ef,
        64'hf1050513_f0c58593,
        64'h44c00613_00003517,
        64'h00003597_80826105,
        64'h45016902_64a200f6,
        64'h10234785_644260e2,
        64'hd7e50805_c763c731,
        64'h8b854105_d59b0107,
        64'h959b93c1_17c20006,
        64'h57839201_16020305,
        64'h061b40c8_00a92023,
        64'h02095913_8d5d1902,
        64'h8d752931_3fff06b7,
        64'h0105151b_f9c7d783,
        64'h00002797_efb50205,
        64'h7793c781_8b89439c,
        64'h93811782_0249079b,
        64'hcb192501_2701dff7,
        64'h77139f21_d007071b,
        64'h777de0bf_f0ef00e7,
        64'h90239381_3ff7071b,
        64'h777d1782_00d71023,
        64'h0329079b_93011702,
        64'h0309071b_00452903,
        64'hc3909381_178227a1,
        64'h842e56fd_415c00e7,
        64'h80234739_938100d7,
        64'h10231782_930192c1,
        64'h02e7879b_170216c2,
        64'h0067871b_eb758b05,
        64'h43189301_17020247,
        64'h871b415c_0ef71263,
        64'h84aa1117_87931111,
        64'h17b70207_ac235158,
        64'h00002797_14050063,
        64'he04ae426_e822ec06,
        64'h11018082_bdf9852e,
        64'hf4f585e3_c0078793,
        64'hf8e58de3_10078713,
        64'hf4f58de3_808283a7,
        64'h8513eee6_8fe381a7,
        64'h85134705_03454683,
        64'h808231b0_05138082,
        64'h61b00513_f0f70ce3,
        64'h63a00513_47850345,
        64'h4703b715_852efcf5,
        64'h8ce38007_8793f8d5,
        64'h8ce34006_8693fee5,
        64'h84e39007_87136789,
        64'hfeb771e3_fee58be3,
        64'h70078713_808203a5,
        64'he513f4f5_9ae35007,
        64'h879300e5_86633007,
        64'h8713b78d_fce587e3,
        64'hd0070713_f6f588e3,
        64'h61a50513_60050793,
        64'h65218082_f6f59fe3,
        64'h20900513_20000793,
        64'hf8f586e3_10200513,
        64'h10000793_808201a5,
        64'he513f8f5_9ee3a007,
        64'h8793fae5_83e39097,
        64'h85139007_87130ab7,
        64'h6f6300e5_8e63b007,
        64'h87138082_fae59fe3,
        64'h90278513_90078713,
        64'hfce586e3_33a78513,
        64'h30078713_fce58ce3,
        64'ha1a78513_a0078713,
        64'h67ad06b7_f66308f5,
        64'h8c637007_07936725,
        64'h0ab77463_04e58f63,
        64'h70068713_668d8082,
        64'h852e12f5_856351b0,
        64'h05135000_079300f5,
        64'h896371a0_05137000,
        64'h07930ef5_8e636000,
        64'h079308b7_f96310f5,
        64'h8e633000_079306b7,
        64'h6c638007_87131207,
        64'h09638005_871b04b7,
        64'h62630ee5_8a632007,
        64'h87136785_80820141,
        64'h45051ce7_a4234705,
        64'h00002797_640260a2,
        64'hcb3ff0ef_1b450513,
        64'h1b058593_0b500613,
        64'h00003517_00003597,
        64'h80820141_45051ee7,
        64'haa234705_00002797,
        64'h640260a2_cdfff0ef,
        64'h1e050513_1dc58593,
        64'h0b400613_00003517,
        64'h00003597_b791472d,
        64'hf406d5e3_47050257,
        64'h9693f406_cae34735,
        64'h02679693_b781dfff,
        64'hf0ef0c80_0513f4e7,
        64'h96e38ff5_40000737,
        64'hc00006b7_541c8082,
        64'h01414505_640260a2,
        64'hb70900f6_002347c1,
        64'h80820141_00e79023,
        64'h20000713_938126d7,
        64'h18231782_00002717,
        64'h46cd0007_10232791,
        64'h93010006_90231702,
        64'h928103a7_871b1682,
        64'h00c71023_3ff6061b,
        64'h0387869b_9301767d,
        64'h170200c6_90230367,
        64'h871b9281_16820347,
        64'h869b6402_60a2405c,
        64'h00e78023_93811782,
        64'h0287879b_4741405c,
        64'h00e78023_93811782,
        64'h0297879b_eff00613,
        64'h405c0a06_d5630277,
        64'h9693473d_541ce941,
        64'h654010ef_8522a805,
        64'h85930006_25b70af7,
        64'h06634789_03644703,
        64'h00f68023_9281d410,
        64'h47bd1682_0296869b,
        64'h43109301_02f40b23,
        64'h0ff7f793_17020406,
        64'h871b0007_d7839381,
        64'h17820fe6_879bffed,
        64'h8b850007_47839301,
        64'h170202f6_871b4054,
        64'h00e78023_93811782,
        64'h02f7879b_4705405c,
        64'hf19ff0ef_3e800513,
        64'h00060023_10e78063,
        64'h92014709_0ff7f793,
        64'h06043823_06042223,
        64'h1602d478_0296061b,
        64'h47190007_d7839381,
        64'h02e40023_17820fe6,
        64'h079b0205_c703cc58,
        64'hcc14c848_01042823,
        64'h01142623_d05cc050,
        64'h00641023_1117879b,
        64'h111117b7_c41c4d94,
        64'h49c80105_a80300c5,
        64'ha8830005_d3034dd8,
        64'h842a459c_1c058c63,
        64'h3c07a223_00002797,
        64'h1a050c63_e022e406,
        64'h11418082_f5450513,
        64'h00002517_8082f825,
        64'h05130000_25178082,
        64'h00e78363_45010247,
        64'hd783f727_87930000,
        64'h279702a7_8163872a,
        64'hf807d783_00002797,
        64'h8082fea7_ebe38f99,
        64'hfda78793_00000797,
        64'h02f50533_02800793,
        64'hfee78ee3_ff86b703,
        64'h0200c6b7_ff87b783,
        64'h0200c7b7_8082ff87,
        64'hb5030200_c7b78082,
        64'h612570a2_a1bff0ef,
        64'he43aecc6_e8c2e4be,
        64'hf40672c5_0513567d,
        64'h080c86b2_1838ec2e,
        64'he0bafc36_fffff517,
        64'he82a711d_a43ff06f,
        64'h72e50513_fffff517,
        64'h85aa862e_86b28736,
        64'h80826105_60e2a5df,
        64'hf0efec06_a6450513,
        64'h002c567d_872e0000,
        64'h051786aa_11018082,
        64'h616160e2_a7bff0ef,
        64'he43ae4c6_e0c2fc3e,
        64'hec061038_77450513,
        64'hf83affff_f51785aa,
        64'h862e86b2_f436715d,
        64'h80826161_60e2aa5f,
        64'hf0efe43a_e4c6e0c2,
        64'hfc3eec06_7a250513,
        64'h1018567d_f83af032,
        64'hfffff517_85aa86ae,
        64'hf436715d_80826125,
        64'h60e2ad1f_f0efe43a,
        64'hecc6e8c2_e4beec06,
        64'hae650513_567d1038,
        64'h858ae0ba_f832f42e,
        64'h00000517_86aafc36,
        64'h711db31d_4809b32d,
        64'h4821bb1d_48410206,
        64'he693bb49_8da29902,
        64'h02500513_85d2866e,
        64'h86ce001d_8413b7d5,
        64'h86222c85_99020016,
        64'h04130200_051385d2,
        64'h86cebb6d_8db28aea,
        64'h018ce563_c019fc08,
        64'h9de3fff8_869bfe0a,
        64'h82e3c519_01b70633,
        64'h00074503_78a27702,
        64'h990285d2_86cef83a,
        64'hf03af446_070588b6,
        64'hb7e178c2_8df28cc2,
        64'h77627e02_78229902,
        64'h02000513_85d286ce,
        64'h866ef072_f442f846,
        64'hfc3a001d_8e13b7c9,
        64'h0785a081_40ed8db3,
        64'h8cc2018c_e863001c,
        64'h881be411_0006841b,
        64'h8a890006_0c9b8666,
        64'h011cf363_8646000a,
        64'h886340e7_8cbb2a81,
        64'h4006fa93_02f61b63,
        64'hc1990007_c58387ba,
        64'h00f70633_93810208,
        64'h97930008_856357fd,
        64'h000ab703_008a8d13,
        64'hb7cd8ca2_2b059902,
        64'h02000513_85d286ce,
        64'h001c8413_8666b559,
        64'h8de68aea_018b6563,
        64'hc0199902_001d8c93,
        64'h008a8d13_85d2866e,
        64'h86ce000a_c503ff87,
        64'h64e3001d_8d130017,
        64'h0b1b8dea_875a9902,
        64'h02000513_85d286ce,
        64'h866ea809_4705e00d,
        64'h4b050006_841b8a89,
        64'hb7ed8f7d_67e2dbe5,
        64'h0807f793_b7699301,
        64'h4781e062_e4361702,
        64'h0ff77713_ca09000a,
        64'ha7030407_f613b755,
        64'he062e436_4781000a,
        64'hb703c719_1007f713,
        64'hbde54781_e062e436,
        64'h000ab703_c719bff1,
        64'h000aa783_b7cd000a,
        64'h9783c781_0807f793,
        64'hbfd940e6_073b93fd,
        64'he062e436_00e7c633,
        64'h41f7d71b_000ac783,
        64'hcf090406_f713b789,
        64'hbb7ff0ef_854a85d2,
        64'h866e86ce_93fd40e6,
        64'h073300f7_463343f7,
        64'hd713e062_e436000a,
        64'hb783c31d_87b61006,
        64'hf713b5dd_07800793,
        64'heef509e3_07500793,
        64'ha89d4841_e03ee436,
        64'h008a8413_000ab703,
        64'h47c10216_e693d4f5,
        64'h1ae30700_0793f0f5,
        64'h0ce306f0_079302a7,
        64'he56312f5_0f630730,
        64'h0793b71d_06400793,
        64'h0ef50663_06300793,
        64'hbddd0c06_e6938082,
        64'h614d6da6_6d466ce6,
        64'h7c067ba6_7b467ae6,
        64'h6a0a69aa_694a64ea,
        64'h000d851b_740a70aa,
        64'h99024501_85d286ce,
        64'hfff98613_013de463,
        64'h866eda05_17e30004,
        64'hc5038aa2_8daacf5f,
        64'hf0ef854a_85d2866e,
        64'h86ce93fd_40e60733,
        64'h00f74633_43f7d713,
        64'he062e436_000ab783,
        64'hcf4510c5_1c630640,
        64'h061300c5_0663008a,
        64'h84130208_58132701,
        64'h87b60690_06131802,
        64'h2006f713_9af9c391,
        64'h4006f793_9acd00f5,
        64'h03630640_079300f5,
        64'h07634829_9abd0690,
        64'h07932ef5_04630620,
        64'h07932ef5_066306f0,
        64'h07932ef5_06630580,
        64'h07932ef5_0c630780,
        64'h0793e4f5_14e30580,
        64'h07932ef5_08630250,
        64'h07930ca7_ef6300f5,
        64'h0c630620_07930ea7,
        64'hec6302f5_02630017,
        64'h04930690_07930007,
        64'h45030806_e6930ef6,
        64'h0e630014_c603a039,
        64'h00248713_3006e693,
        64'ha8211006_e69300f6,
        64'h05630014_c603b7e9,
        64'h07a00613_00c78963,
        64'h07400613_bf6584ba,
        64'hbf758abe_04892881,
        64'h48810008_d363008a,
        64'h8793000a_a88300f6,
        64'h1d6302a0_0793a899,
        64'h872604c7_806306a0,
        64'h061304c7_8c630680,
        64'h061302f6_6d6304c7,
        64'h86630014_871306c0,
        64'h06130004_c783fef6,
        64'h71e30ff7_f793fd07,
        64'h079b0014_85930004,
        64'hc70300e8_88bbfd08,
        64'h889b84ae_031b88bb,
        64'hb77584b2_8aba40f0,
        64'h0c3b0026_e6930007,
        64'hd6630007_8c1b008a,
        64'h8713000a_a783fce7,
        64'h96e34c01_02a00713,
        64'ha8254625_84ba06f5,
        64'hee634006_e6930ff7,
        64'hf793fd06_079b0014,
        64'h871345a5_0014c603,
        64'h06f71763_488102e0,
        64'h07930004_c703fef6,
        64'h71e30ff7_f793fd07,
        64'h079b0014_85930004,
        64'hc70300e3_0c3bfd03,
        64'h031b84ae_038b833b,
        64'hbf750106_e693b7c9,
        64'h0086e693_b7e10046,
        64'he693b7f9_0026e693,
        64'ha0254625_4c0106e5,
        64'he96345a5_0ff77713,
        64'hfd07871b_02a78563,
        64'h02b78463_fcf76fe3,
        64'h02e78563_00148613,
        64'h0004c783_84b20016,
        64'he6930287_91630300,
        64'h04130287_8f6302d0,
        64'h0413a821_02300513,
        64'h02000593_02b00713,
        64'h4681a155_85d2866e,
        64'h86ce001d_841300f5,
        64'h08630485_02500793,
        64'hac814ba9_ec3e4d81,
        64'hfffb0793_6b41cc89,
        64'h09130000_0917e589,
        64'h892a8aba_84b689b2,
        64'h8a2ee4ee_e8eaece6,
        64'hf0e2f4de_f8daf122,
        64'hf506fcd6_e152e54e,
        64'he94aed26_71718082,
        64'h9c7ff06f_c119b7e1,
        64'h006e033b_80826161,
        64'h60a6d17f_f0ef887e,
        64'h10180008_089be43a,
        64'he876e046_4746fc57,
        64'h9de3c319_fe6f0fa3,
        64'h9f3e0ff3_73130201,
        64'h0f130785_03075733,
        64'h0303031b_03e3ee63,
        64'h0fff7313_03077f33,
        64'h02000293_ff630e1b,
        64'h43a54781_04100313,
        64'h000e0463_06100313,
        64'h020efe13_c7214781,
        64'h00030463_400ef313,
        64'hfefefe93_e3194ee6,
        64'h8fbee486_715db7e1,
        64'h006e033b_80826161,
        64'h60a6d97f_f0ef887e,
        64'h10180008_089be43a,
        64'he876e046_4746fc57,
        64'h9de3c319_fe6f0fa3,
        64'h9f3e0ff3_73130201,
        64'h0f130785_03075733,
        64'h0303031b_03e3ee63,
        64'h0fff7313_03077f33,
        64'h02000293_ff630e1b,
        64'h43a54781_04100313,
        64'h000e0463_06100313,
        64'h020efe13_c7214781,
        64'h00030463_400ef313,
        64'hfefefe93_e3194ee6,
        64'h8fbee486_715db7a9,
        64'h86229b02_00160413,
        64'h02000513_85de86e2,
        64'hb7919b02_85de86e2,
        64'h00094503_b7ed4154,
        64'h0cb30209_59130209,
        64'h9913bf89_ff27e3e3,
        64'h009c87b3_84ea0014,
        64'h8d136722_9b02e43a,
        64'h02000513_85de86e2,
        64'h8626b7ad_00d60023,
        64'h00870633_da3d0087,
        64'hf613bf9d_02b00613,
        64'h008706b3_c6110047,
        64'hf613bfa1_06200613,
        64'h008706b3_f886ece3,
        64'h46fdf6d8_98e34689,
        64'hb7bd0580_06130087,
        64'h06b3fa86_e7e346fd,
        64'h80826165_85326d42,
        64'h6ce27c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a60b37,
        64'he1634156_07b30209,
        64'hd9931982_000a0963,
        64'h00940633_0b2c9663,
        64'h197d412d_06330124,
        64'h8d33fff7_0c930087,
        64'h0933cbcd_84d68b8d,
        64'h040500c6_802302d0,
        64'h06130087_06b30808,
        64'h046300d4_0b630200,
        64'h06930405_00c68023,
        64'h03000613_008706b3,
        64'h0286e663_46fd0405,
        64'h00c68023_07800613,
        64'h008706b3_0486e063,
        64'h46fdead1_0207f693,
        64'h0ad89663_46c14401,
        64'hbf55fe6e_0fa30087,
        64'h0e330405_a0e902c8,
        64'h9a638436_460902c8,
        64'h81631479_4641c285,
        64'hfff40693_02869563,
        64'h92810209_96930086,
        64'h87639281_1682cc0d,
        64'hee154007_f613ca3d,
        64'h0107f613_02b41e63,
        64'h00a47463_c6090300,
        64'h03130200_05939101,
        64'h02099513_fea469e3,
        64'hfe6e0fa3_00870e33,
        64'h040500b4_0963a801,
        64'h03000313_02000593,
        64'h91010206_951339fd,
        64'hc19100c7_f5930008,
        64'h1563c619_00098963,
        64'h0017f613_040a1a63,
        64'h59e656c6_8ab28bae,
        64'h8b2a8c36_2a01e86a,
        64'hec66e8ca_eca6f486,
        64'hf062f45e_f85afc56,
        64'h0027fa13_e4cee0d2,
        64'h478a843e_f0a27159,
        64'h80828302_658c0005,
        64'hb303c509_80828082,
        64'h00a58023_95b200d6,
        64'h7563bbe1_02f000ef,
        64'hd1850513_00004517,
        64'hbd35adc5_051385a6,
        64'h00004517_047000ef,
        64'had050513_00004517,
        64'hcd0984aa_dd1ff0ef,
        64'h8552865a_020aa583,
        64'h063000ef_d3450513,
        64'h00004517_f57990e3,
        64'h08048493_077000ef,
        64'h2985b325_05130000,
        64'h4517ff2c_17e30890,
        64'h00ef0905_cd450513,
        64'h00004517_00094583,
        64'h07048c13_02848913,
        64'h0a3000ef_d5c50513,
        64'h00004517_0af000ef,
        64'hd5050513_00004517,
        64'h708c0bd0_00efd465,
        64'h05130000_45176c8c,
        64'h0cb000ef_d3c50513,
        64'h00004517_688cff2c,
        64'h17e30dd0_00ef0905,
        64'hd2850513_00004517,
        64'h00094583_01090c13,
        64'h0f3000ef_d4450513,
        64'h00004517_fe9917e3,
        64'h103000ef_0905d4e5,
        64'h05130000_45170009,
        64'h4583ff04_89131190,
        64'h00efd425_05130000,
        64'h45171250_00efd385,
        64'h051385ce_00004517,
        64'hbf15d245_051385ce,
        64'h00004517_13f000ef,
        64'hbc850513_00004517,
        64'hcd094b91_080489aa,
        64'h8a8aecff_f0ef850a,
        64'h46057101_44ac1610,
        64'h00efd325_05130000,
        64'h451745d6_16f000ef,
        64'hd2050513_00004517,
        64'h45c617d0_00efd065,
        64'h05130000_451765a6,
        64'h18b000ef_cfc50513,
        64'h00004517_75821990,
        64'h00efcf25_05130000,
        64'h451765e2_1a7000ef,
        64'hce850513_00004517,
        64'h45d21b50_00efcde5,
        64'h05130000_451745c2,
        64'h1c3000ef_cd450513,
        64'h00004517_45b21d10,
        64'h00efcca5_05130000,
        64'h451745a2_1df000ef,
        64'hcc050513_00004517,
        64'h65821ed0_00efcae5,
        64'h05130000_4517b755,
        64'h54f91fd0_00efc9e5,
        64'h05130000_4517fa84,
        64'h358320d0_00efc965,
        64'h05130000_4517faa4,
        64'h3423c11d_f99ff0ef,
        64'h848a850a_45854605,
        64'h710122d0_00efc9e5,
        64'h05130000_45178082,
        64'h61256c42_6be27b02,
        64'h7aa27a42_79e26906,
        64'h64a66446_852660e6,
        64'hfa040113_54fd2590,
        64'h00efca25_05130000,
        64'h4517c51d_f73ff0ef,
        64'h8b2e8a2a_1080e862,
        64'hec5ef456_fc4ee0ca,
        64'he4a6ec86_f05af852,
        64'he8a2711d_80824501,
        64'hbfc94501_28f000ef,
        64'hcb850513_00004517,
        64'hb7cd5575_29f000ef,
        64'hca850513_00004517,
        64'hc9091260_10ef8522,
        64'h80820141_640260a2,
        64'h55792bd0_00efcae5,
        64'h05130000_4517cd01,
        64'h41b000ef_8522c704,
        64'h041341d0_00003417,
        64'hc18d557d_85aa3fb0,
        64'h00ef4501_2e7000ef,
        64'he022e406_cc650513,
        64'h11410000_45178082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_00a78223,
        64'h0ff57513_00d78023,
        64'h0085551b_0ff57693,
        64'h00d78623_f8000693,
        64'h00078223_01e71793,
        64'h470d02b5_553b0045,
        64'h959b8082_00a78023,
        64'hdf650207_77130147,
        64'hc70307fa_478d8082,
        64'h02057513_0147c503,
        64'h07fa478d_80820005,
        64'h45038082_00b50023,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_100004b7,
        64'h18858593_00003597,
        64'hf1402573_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_3ad020ef,
        64'h40000137_03249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
