/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 3532;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_00000001,
        64'h05f5e100_e0101000,
        64'h00000001_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000001_05f5e100,
        64'he0100000_00000000,
        64'h00000030_00003000,
        64'h00000020_00002000,
        64'h00000010_00001000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_322d746c,
        64'h75616665_642d6972,
        64'h742c786e_6c780074,
        64'h6c756166_65642d69,
        64'h72742c78_6e6c7800,
        64'h6c617564_2d73692c,
        64'h786e6c78_00746e65,
        64'h73657270_2d747075,
        64'h72726574_6e692c78,
        64'h6e6c7800_68746469,
        64'h772d326f_6970672c,
        64'h786e6c78_00687464,
        64'h69772d6f_6970672c,
        64'h786e6c78_00322d74,
        64'h6c756166_65642d74,
        64'h756f642c_786e6c78,
        64'h00746c75_61666564,
        64'h2d74756f_642c786e,
        64'h6c780032_2d737475,
        64'h706e692d_6c6c612c,
        64'h786e6c78_00737475,
        64'h706e692d_6c6c612c,
        64'h786e6c78_0072656c,
        64'h6c6f7274_6e6f632d,
        64'h6f697067_00736c6c,
        64'h65632d6f_69706723,
        64'h0070772d_656c6261,
        64'h73696400_7365676e,
        64'h61722d65_6761746c,
        64'h6f760079_636e6575,
        64'h71657266_2d78616d,
        64'h2d697073_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_5a020000,
        64'h04000000_03000000,
        64'hffffffff_49020000,
        64'h04000000_03000000,
        64'h01000000_3c020000,
        64'h04000000_03000000,
        64'h00000000_25020000,
        64'h04000000_03000000,
        64'h08000000_14020000,
        64'h04000000_03000000,
        64'h08000000_04020000,
        64'h04000000_03000000,
        64'h00000000_f0010000,
        64'h04000000_03000000,
        64'h00000000_de010000,
        64'h04000000_03000000,
        64'h00000000_cc010000,
        64'h04000000_03000000,
        64'h00000000_bc010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h000000c1_00000000,
        64'h67000000_10000000,
        64'h03000000_ac010000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'ha0010000_04000000,
        64'h03000000_00000030,
        64'h30303030_30316340,
        64'h6f697067_01000000,
        64'h02000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_03000000,
        64'h52010000_04000000,
        64'h03000000_00000000,
        64'h64656c62_61736964,
        64'h6b000000_09000000,
        64'h03000000_00100000,
        64'h00000000_00b000e0,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00006d65_672c736e,
        64'h6463006d_65672d71,
        64'h6e797a2c_736e6463,
        64'h1b000000_17000000,
        64'h03000000_00000030,
        64'h30306230_30306540,
        64'h74656e72_65687465,
        64'h01000000_02000000,
        64'h02000000_95010000,
        64'h00000000_03000000,
        64'he40c0000_e40c0000,
        64'h86010000_08000000,
        64'h03000000_20bcbe00,
        64'h74010000_04000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00000000,
        64'h746f6c73_2d697073,
        64'h2d636d6d_1b000000,
        64'h0d000000_03000000,
        64'h00000030_40636d6d,
        64'h01000000_00100000,
        64'h00000000_000010e0,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_52010000,
        64'h04000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h00000000_64656c62,
        64'h61736964_6b000000,
        64'h09000000_03000000,
        64'h00000061_392e382d,
        64'h69636864_732c6e61,
        64'h73617261_1b000000,
        64'h12000000_03000000,
        64'h00000000_30303030,
        64'h30313065_40636d6d,
        64'h01000000_02000000,
        64'h00100000_00000000,
        64'h00d000e0_00000000,
        64'h67000000_10000000,
        64'h03000000_02000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h64656c62_61736964,
        64'h6b000000_09000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_0000302e,
        64'h312d6970_73712d71,
        64'h6e797a2c_786e6c78,
        64'h1b000000_13000000,
        64'h03000000_00000000,
        64'h30303064_30303065,
        64'h40697073_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_005a6202,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_000000c0,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30306340,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000030_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h31407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_005a6202,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'hc0e1e400_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30634074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h08090000_6d020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h40090000_38000000,
        64'had0b0000_edfe0dd0,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_6e6f6974,
        64'h706f5f73_70647378,
        64'h000a6425_202c7325,
        64'h203a7472_65737341,
        64'h00632e73_70647378,
        64'hffffb41e_ffffbaba,
        64'hffffbaba_ffffb41e,
        64'hffffbaba_ffffb8a4,
        64'hffffbaba_ffffbaba,
        64'hffffb9de_ffffb41e,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffb41e,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffb41e_ffffb7e0,
        64'hffffb41e_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffb41e_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffbaba,
        64'hffffbaba_ffffba8e,
        64'hffffb408_ffffb420,
        64'hffffb420_ffffb420,
        64'hffffb420_ffffb420,
        64'hffffb3d8_ffffb420,
        64'hffffb420_ffffb420,
        64'hffffb420_ffffb420,
        64'hffffb420_ffffb420,
        64'hffffb358_ffffb420,
        64'hffffb3f0_ffffb420,
        64'hffffb398_ffffb1a4,
        64'hffffb23a_ffffb23a,
        64'hffffb1c2_ffffb23a,
        64'hffffb1e0_ffffb23a,
        64'hffffb23a_ffffb23a,
        64'hffffb23a_ffffb23a,
        64'hffffb23a_ffffb23a,
        64'hffffb21c_ffffb23a,
        64'hffffb23a_ffffb1fe,
        64'h00000a21_656e6f44,
        64'h00000a2e_2e2e6567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f43,
        64'h00000000_00000000,
        64'h20202020_20202020,
        64'h203a656d_616e090a,
        64'h00586c6c_36313025,
        64'h2020203a_73657475,
        64'h62697274_7461090a,
        64'h00000000_00007525,
        64'h20202020_203a6162,
        64'h6c207473_616c090a,
        64'h00000000_00007525,
        64'h20202020_3a61626c,
        64'h20747372_6966090a,
        64'h00000000_00002020,
        64'h20202020_2020203a,
        64'h64697567_206e6f69,
        64'h74697472_6170090a,
        64'h00000000_58323025,
        64'h00000000_00002020,
        64'h20203a64_69756720,
        64'h65707974_206e6f69,
        64'h74697472_6170090a,
        64'h00006425_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h7825203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h000a5838_25202020,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702065_7a697309,
        64'h000a5838_25203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20726562_6d756e09,
        64'h00000000_000a586c,
        64'h6c363130_25202020,
        64'h203a6162_6c207365,
        64'h6972746e_65206e6f,
        64'h69746974_72617009,
        64'h00000000_0a756c6c,
        64'h25202020_3a61646c,
        64'h2070756b_63616209,
        64'h00000000_0a756c6c,
        64'h2520203a_61626c20,
        64'h746e6572_72756309,
        64'h00000000_0a583830,
        64'h25202020_20203a64,
        64'h65767265_73657209,
        64'h00000000_0a583830,
        64'h25202020_3a726564,
        64'h6165685f_63726309,
        64'h00000000_0a583830,
        64'h25202020_20202020,
        64'h20203a65_7a697309,
        64'h00000000_0a583830,
        64'h25202020_20203a6e,
        64'h6f697369_76657209,
        64'h00000000_0000000a,
        64'h00000000_00006325,
        64'h00202020_203a6572,
        64'h7574616e_67697309,
        64'h00000000_0a3a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20545047,
        64'h00000000_0000000a,
        64'h6425203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_635f6473,
        64'h00000000_00000000,
        64'h0a216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_00000000,
        64'h0a216465_7a696c61,
        64'h6974696e_69204453,
        64'h00000000_000a676e,
        64'h69746978_65202e2e,
        64'h2e445320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f43,
        64'h00000000_0a642520,
        64'h3a737574_61747320,
        64'h2c64656c_69616620,
        64'h64616552_20304453,
        64'h00000000_0a216465,
        64'h65636375_73206e6f,
        64'h6974617a_696c6169,
        64'h74696e49_20304453,
        64'h00000000_000a6425,
        64'h203a7375_74617473,
        64'h202c6465_6c696166,
        64'h206e6f69_74617a69,
        64'h6c616974_696e6920,
        64'h64726163_20304453,
        64'h0000000a_6425203a,
        64'h73757461_7473202c,
        64'h64656c69_6166206c,
        64'h61697469_6e692067,
        64'h69666e6f_63204453,
        64'h00000000_0000000a,
        64'h2164656c_69616620,
        64'h6769666e_6f632070,
        64'h756b6f6f_6c204453,
        64'h00000000_000a2e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e49,
        64'h00000000_0000000a,
        64'h6c696166_20746f6f,
        64'h62206567_61747320,
        64'h6f72657a_20514e59,
        64'h5a20656e_61697241,
        64'h00000020_58323025,
        64'h00000000_0000000a,
        64'h786c6c25_78304045,
        64'h5341425f_4d415244,
        64'h00000000_0000000a,
        64'h000a6425_202c6425,
        64'h00000000_002e2e2e,
        64'h00000000_00000a72,
        64'h6564616f_6c746f6f,
        64'h42206567_61745320,
        64'h6f72655a_20514e59,
        64'h5a20656e_61697241,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623a14f,
        64'hc0ef4505_a031fef4,
        64'h26234785_e7892781,
        64'h0807f793_278187aa,
        64'haa5fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'h0001a011_f6e7fee3,
        64'h02700793_0ff7f713,
        64'hfe944783_fef404a3,
        64'h2785fe94_4783cf99,
        64'h27810407_f7932781,
        64'h87aaadff_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h3783a0ad_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hae5fd0ef_fd843503,
        64'h50078593_67854601,
        64'h4685a829_fef42623,
        64'h87aaafff_d0effd84,
        64'h35033007_85936785,
        64'h46014685_00f71f63,
        64'h4785873e_0347c783,
        64'hfd843783_a8adfe04,
        64'h04a3ad0f_c0ef4505,
        64'hb87fe0ef_853e03e0,
        64'h0593863a_fe645703,
        64'h43dcfd84_3783fef4,
        64'h13230407_e793fe64,
        64'h5783fef4_132387aa,
        64'hb75fe0ef_853e03e0,
        64'h059343dc_fd843783,
        64'hc2e19423_4741bc5f,
        64'he0ef853e_4591863a,
        64'hfea45703_43dcfd84,
        64'h3783fef4_15238ff9,
        64'h17fd6785_fea45703,
        64'hfef41523_0017979b,
        64'hfea45783_aa254785,
        64'hc2e1a223_470593af,
        64'hc0ef78a5_05130000,
        64'h05177825_85930000,
        64'h05974b60_0613a015,
        64'h02f71a63_478d873e,
        64'h0377c783_fd843783,
        64'hfef41523_04000793,
        64'hc201a223_aaa54785,
        64'hc2e1a223_470597af,
        64'hc0ef7ca5_05130000,
        64'h05177c25_85930000,
        64'h05974b50_0613a015,
        64'h04f71363_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_c201a223,
        64'hcf91fd84_3783fca4,
        64'h3c231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_beffe0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fd843783,
        64'hcaffe0ef_853e0300,
        64'h05934609_43dcfd84,
        64'h3783dfc5_27818b89,
        64'hfe842783_a83dfef4,
        64'h26234785_cd3fe0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c385_27818ff9,
        64'h67a1fe84_2703fef4,
        64'h242387aa_cc1fe0ef,
        64'h853e0300_059343dc,
        64'hfd843783_a8bdfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aacc7f_d0effd84,
        64'h35036000_0593863e,
        64'h4681fd44_2783fcf4,
        64'h2a2387ae_fca43c23,
        64'h1800f022_f4067179,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aacb5f_e0ef853e,
        64'h93811782_278127c1,
        64'h43dcfc84_3783d75f,
        64'he0ef853e_03000593,
        64'h460943dc_fc843783,
        64'hdfc52781_8b89fdc4,
        64'h2783a83d_fef42623,
        64'h4785d99f_e0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fc843783,
        64'hc3852781_8ff967a1,
        64'hfdc42703_fcf42e23,
        64'h87aad87f_e0ef853e,
        64'h03000593_43dcfc84,
        64'h3783a8bd_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hd8dfd0ef_fc843503,
        64'h80078593_6785863e,
        64'h4685fe44_2783c2e1,
        64'h94234745_7010d073,
        64'h70105073_0ff0000f,
        64'hfc2fe0ef_fc843503,
        64'h85befc04_36032781,
        64'hfe245783_e23fe0ef,
        64'h853e4591_863afe04,
        64'h570343dc_fc843783,
        64'hfef41023_8ff917fd,
        64'h6785fe04_5703fef4,
        64'h10232000_0793fef4,
        64'h11234785_fce7dee3,
        64'h1ff00793_0007871b,
        64'hfe842783_fef42423,
        64'h2785fe84_27830007,
        64'h802397ba_fc043703,
        64'hfe842783_a2354785,
        64'hc2e1a223_4705bc2f,
        64'hc0efa125_05130000,
        64'h1517a0a5_85930000,
        64'h15973750_0613a835,
        64'hfe042423_c201a223,
        64'haaa14785_c2e1a223,
        64'h4705beef_c0efa3e5,
        64'h05130000_1517a365,
        64'h85930000_15973740,
        64'h0613a015_02f71963,
        64'h11178793_111117b7,
        64'h873e53dc_fc843783,
        64'hc201a223_cf91fc84,
        64'h3783fe04_2223fcb4,
        64'h3023fca4_34230080,
        64'hf822fc06_71398082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'ha019fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaecbf,
        64'hd0effd84_3503a007,
        64'h859367ad_46014681,
        64'ha03dfef4_26234785,
        64'ha82d4785_c2e1a223,
        64'h4705c86f_c0efad65,
        64'h05130000_1517ace5,
        64'h85930000_15973450,
        64'h0613a015_c79d2781,
        64'hfec42783_fef42623,
        64'h87aaf17f_d0effd84,
        64'h35037007_8593678d,
        64'h863e4681_4bbcfd84,
        64'h3783c201_a223a061,
        64'h4785c2e1_a2234705,
        64'hcd4fc0ef_b2450513,
        64'h00001517_b1c58593,
        64'h00001597_34400613,
        64'ha01504f7_1a631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783c201,
        64'ha223cf91_fd843783,
        64'hfca43c23_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_853efe84,
        64'h2783fe04_2423fedf,
        64'he0ef853a_02c00593,
        64'h863e93c1_17c20047,
        64'he793fe44_578343d8,
        64'hfd843783_fef41223,
        64'h87aafd7f_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783d3e5_27818b89,
        64'h2781fe64_5783fef4,
        64'h132387aa_ff9fe0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_a821fef4,
        64'h132387aa_810ff0ef,
        64'h853e02c0_059343dc,
        64'hfd843783_85aff0ef,
        64'h853e02c0_0593863a,
        64'hfe445703_43dcfd84,
        64'h3783fef4_12230017,
        64'he79393c1_17c28fd9,
        64'hfe445783_fec45703,
        64'hfef41623_f007f793,
        64'hfec45783_fef41623,
        64'h0087979b_fec45783,
        64'hfef41223_0ff7f793,
        64'hfe445783_fef41223,
        64'h87aa876f_f0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783a0a5_8c2ff0ef,
        64'h853e02c0_0593863a,
        64'hfe445703_43dcfd84,
        64'h3783fef4_12230017,
        64'he79393c1_17c28fd9,
        64'hfe445783_93410307,
        64'h97138fd9_fe245783,
        64'hfec45703_fef41623,
        64'hf007f793_fec45783,
        64'hfef41623_0087979b,
        64'hfec45783_fef41123,
        64'h0c07f793_fe245783,
        64'hfef41123_0067979b,
        64'hfe245783_fef41123,
        64'h0087d79b_fec45783,
        64'hfef41223_03f7f793,
        64'hfe445783_fef41223,
        64'h87aa90ef_f0ef853e,
        64'h02c00593_43dcfd84,
        64'h378308f7_1e634789,
        64'h873e0367_c783fd84,
        64'h3783a249_fef42423,
        64'h478500e7_f6631000,
        64'h07930007_871bfee4,
        64'h5783fae7_fee31000,
        64'h07930007_871bfee4,
        64'h5783fef4_17230017,
        64'h979bfee4_5783a839,
        64'hfef41623_0017d79b,
        64'hfee45783_00e7e963,
        64'h2781fd44_27830007,
        64'h871b02f7_57bb2781,
        64'hfee45783_4798fd84,
        64'h3783a82d_fef41723,
        64'h4785a2ed_fef42423,
        64'h478506e7_fa637fe0,
        64'h07930007_871bfee4,
        64'h5783fae7_ffe37fe0,
        64'h07930007_871bfee4,
        64'h5783fef4_17232785,
        64'hfee45783_a831fef4,
        64'h16230017_d79bfee4,
        64'h578300e7_e9632781,
        64'hfd442783_0007871b,
        64'h02f757bb_2781fee4,
        64'h57834798_fd843783,
        64'ha825fef4_17234785,
        64'hac914785_c2e1a223,
        64'h4705f7ef_c0efdce5,
        64'h05130000_1517dc65,
        64'h85930000_15972d00,
        64'h0613a015_08f71763,
        64'h4789873e_0367c783,
        64'hfd843783_a6aff0ef,
        64'h853e02c0_0593863a,
        64'hfe445703_43dcfd84,
        64'h3783fef4_12239be9,
        64'hfe445783_fef41223,
        64'h87aaa56f_f0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783c201_a223a4c9,
        64'h4785c2e1_a2234705,
        64'hfecfc0ef_e3c50513,
        64'h00001517_e3458593,
        64'h00001597_2cf00613,
        64'ha01506f7_1a631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783c201,
        64'ha223cf91_fd843783,
        64'hfe041623_fcf42a23,
        64'h87aefca4_3c231800,
        64'hf022f406_71798082,
        64'h61657406_70a6853e,
        64'hfec42783_fe042623,
        64'hfef42623_278187aa,
        64'ha6aff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hf9843783_baaff0ef,
        64'h853e0280_0593863a,
        64'h0ff77713_fe442703,
        64'h43dcf984_3783fef4,
        64'h22230047_e793fe44,
        64'h2783fef4_222387aa,
        64'hb9cff0ef_853e0280,
        64'h059343dc_f9843783,
        64'hab7fc0ef_3e800513,
        64'ha09dfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa7080,
        64'h00eff984_350302f7,
        64'h1163479d_873e57fc,
        64'hf9843783_a849fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa0b80_00eff984,
        64'h350385be_5f9cf984,
        64'h3783bc0f_f0ef853e,
        64'h03000593_460943dc,
        64'hf9843783_dfc52781,
        64'h8b89fe44_2783a8d1,
        64'hfef42623_4785be4f,
        64'hf0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hf9843783_c3852781,
        64'h8ff967a1_fe442703,
        64'hfef42223_87aabd2f,
        64'hf0ef853e_03000593,
        64'h43dcf984_3783aa11,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_bd8fe0ef,
        64'hf9843503_60000593,
        64'h863e4681_fe842783,
        64'hdf985007_071b0319,
        64'h7737f984_3783fef4,
        64'h24231007_879b03b9,
        64'h07b7a831_df985007,
        64'h071b0319_7737f984,
        64'h3783fef4_24231007,
        64'h879b03b9_07b702f7,
        64'h10634791_873e57fc,
        64'hf9843783_a099df98,
        64'h2007071b_0bebc737,
        64'hf9843783_fef42423,
        64'h2007879b_03b907b7,
        64'h02f71063_479d873e,
        64'h57fcf984_3783a275,
        64'hfef42623_47851407,
        64'h89632781_fec42783,
        64'hfef42623_87aa1d40,
        64'h00eff984_35035007,
        64'h85930319_77b7df98,
        64'h5007071b_03197737,
        64'hf9843783_ceaff0ef,
        64'h853e0300_05934609,
        64'h43dcf984_3783dfc5,
        64'h27818b89_fe442783,
        64'haafdfef4_26234785,
        64'hd0eff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8f984_3783c385,
        64'h27818ff9_67a1fe44,
        64'h2703fef4_222387aa,
        64'hcfcff0ef_853e0300,
        64'h059343dc_f9843783,
        64'hac3dfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aad02f,
        64'he0eff984_35036000,
        64'h0593863e_4681fe84,
        64'h2783fef4_24231007,
        64'h879b03b9_07b70cf7,
        64'h16634789_873e0347,
        64'hc783f984_3783a451,
        64'hfef42623_47852207,
        64'h85632781_fec42783,
        64'hfef42623_87aa2ac0,
        64'h00eff984_350385be,
        64'h5f9cf984_3783df98,
        64'h0807071b_02faf737,
        64'hf9843783_dc2ff0ef,
        64'h853e0300_05934609,
        64'h43dcf984_3783dfc5,
        64'h27818b89_fe442783,
        64'hacd9fef4_26234785,
        64'hde6ff0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8f984_3783c385,
        64'h27818ff9_67a1fe44,
        64'h2703fef4_222387aa,
        64'hdd4ff0ef_853e0300,
        64'h059343dc_f9843783,
        64'hae19fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aaddaf,
        64'he0eff984_35036000,
        64'h0593863e_4685fe84,
        64'h2783fef4_242337c5,
        64'h810007b7_c2e19423,
        64'h47457010_d0737010,
        64'h50730ff0_000f818f,
        64'hf0eff984_350385be,
        64'h863afa04_07132781,
        64'hfe245783_e7aff0ef,
        64'h853e4591_863afe04,
        64'h570343dc_f9843783,
        64'hfef41023_8ff917fd,
        64'h6785fe04_5703fef4,
        64'h10230400_0793fef4,
        64'h11234785_a65d4785,
        64'hc2e1a223_4705bf3f,
        64'hc0ef2425_05130000,
        64'h151723a5_85930000,
        64'h15972040_0613a015,
        64'h14f71363_4785873e,
        64'h0347c783_f9843783,
        64'hc201a223_aef94785,
        64'hc2e1a223_4705c2bf,
        64'hc0ef27a5_05130000,
        64'h15172725_85930000,
        64'h15972030_0613a015,
        64'h02f71f63_11178793,
        64'h111117b7_873e53dc,
        64'hf9843783_c201a223,
        64'hcf91f984_3783fc04,
        64'h3c23fc04_3823fc04,
        64'h3423fc04_3023fa04,
        64'h3c23fa04_3823fa04,
        64'h3423fa04_3023f8a4,
        64'h3c231880_f0a2f486,
        64'h71598082_61217442,
        64'h70e2853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_ebeff0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fc843783,
        64'hf7eff0ef_853e0300,
        64'h05934609_43dcfc84,
        64'h3783dfc5_27818b89,
        64'hfdc42783_a83dfef4,
        64'h26234785_fa2ff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fc84,
        64'h3783c385_27818ff9,
        64'h67a1fdc4_2703fcf4,
        64'h2e2387aa_f90ff0ef,
        64'h853e0300_059343dc,
        64'hfc843783_a8bdfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaf96f_e0effc84,
        64'h35036000_0593863e,
        64'h4685fe04_27837010,
        64'hd0737010_50730ff0,
        64'h000ffef4_202337c1,
        64'h010007b7_c2e19423,
        64'h47459d4f_f0effc84,
        64'h350385be_fc043603,
        64'h2781fe64_5783835f,
        64'hf0ef853e_4591863a,
        64'hfe445703_43dcfc84,
        64'h3783fef4_12238ff9,
        64'h17fd6785_fe445703,
        64'hfef41223_04000793,
        64'hfef41323_4785fce7,
        64'hdee303f0_07930007,
        64'h871bfe84_2783fef4,
        64'h24232785_fe842783,
        64'h00078023_97bafc04,
        64'h3703fe84_2783aa15,
        64'h4785c2e1_a2234705,
        64'hdd5fc0ef_42450513,
        64'h00001517_41c58593,
        64'h00001597_1a800613,
        64'ha835fe04_2423c201,
        64'ha223a285_4785c2e1,
        64'ha2234705_e01fc0ef,
        64'h45050513_00001517,
        64'h44858593_00001597,
        64'h1a700613_a01502f7,
        64'h19631117_87931111,
        64'h17b7873e_53dcfc84,
        64'h3783c201_a223cf91,
        64'hfc843783_fcb43023,
        64'hfca43423_0080f822,
        64'hfc067139_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623fef4,
        64'h26232781_87aa879f,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfd84,
        64'h3783939f_f0ef853e,
        64'h03e00593_863a9341,
        64'h1742fe84_270343dc,
        64'hfd843783_fef42423,
        64'h8fd9fe84_278357f8,
        64'hfd843783_fef42423,
        64'h8ff917e1_67c1fe84,
        64'h2703fef4_242387aa,
        64'h93dff0ef_853e03e0,
        64'h059343dc_fd843783,
        64'h04f71963_4791873e,
        64'h57fcfd84_3783a15f,
        64'hf0ef853e_02800593,
        64'h863a0ff7_7713fe84,
        64'h270343dc_fd843783,
        64'hfef42423_0027e793,
        64'hfe842783_a039fef4,
        64'h24230207_e793fe84,
        64'h278300f7_1963478d,
        64'h873e0377_c783fd84,
        64'h3783fef4_242387aa,
        64'ha25ff0ef_853e0280,
        64'h059343dc_fd843783,
        64'h93efd0ef_3e800513,
        64'h9f7ff0ef_853e0300,
        64'h05934609_43dcfd84,
        64'h3783dfc5_27818b89,
        64'hfe842783_a8f5fef4,
        64'h26234785_a1bff0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c385_27818ff9,
        64'h67a1fe84_2703fef4,
        64'h242387aa_a09ff0ef,
        64'h853e0300_059343dc,
        64'hfd843783_aa35fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaa0ff_e0effd84,
        64'h35036000_0593863e,
        64'h4681fe44_2783fef4,
        64'h22231007_879b03b7,
        64'h07b7a039_fef42223,
        64'h5007879b_03b707b7,
        64'h00f71963_4791873e,
        64'h57fcfd84_3783a02d,
        64'hfef42223_2007879b,
        64'h03b707b7_a825fef4,
        64'h22236007_879b03b7,
        64'h07b700f7_19634791,
        64'h873e57fc_fd843783,
        64'h02f71763_478d873e,
        64'h0377c783_fd843783,
        64'h02e78ba3_4709fd84,
        64'h3783a031_02e78ba3,
        64'h470dfd84_378300f7,
        64'h186347a1_873e4bdc,
        64'hfd843783_00f71f63,
        64'h4795873e_0347c783,
        64'hfd843783_02f71763,
        64'h4789873e_0367c783,
        64'hfd843783_a431fef4,
        64'h26234785_12078c63,
        64'h2781fec4_2783fef4,
        64'h262387aa_ae1fe0ef,
        64'hfd843503_60078593,
        64'h67a1863e_4681fe44,
        64'h2783fef4_22230377,
        64'hc783fd84_378302e7,
        64'h8ba34709_fd843783,
        64'hac81fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aab23f,
        64'he0effd84_35037007,
        64'h8593678d_863e4681,
        64'h4bbcfd84_378306f7,
        64'h1b634785_873e0347,
        64'hc783fd84_3783a479,
        64'hfe042623_00e7e563,
        64'h478d873e_4bdcfd84,
        64'h3783a45d_4785c2e1,
        64'ha2234705_900fd0ef,
        64'h75050513_00001517,
        64'h74858593_00001597,
        64'h11b00613_a01502f7,
        64'h1e634789_873e0367,
        64'hc783fd84_3783c201,
        64'ha223acf9_4785c2e1,
        64'ha2234705_938fd0ef,
        64'h78850513_00001517,
        64'h78058593_00001597,
        64'h11a00613_a01502f7,
        64'h1f631117_87931111,
        64'h17b7873e_53dcfd84,
        64'h3783c201_a223cf91,
        64'hfd843783_fca43c23,
        64'h1800f022_f4067179,
        64'h80826145_740270a2,
        64'h853efec4_2783fe04,
        64'h2623fef4_26232781,
        64'h87aabadf_f0ef853e,
        64'h93811782_278127c1,
        64'h43dcfd84_3783c6df,
        64'hf0ef853e_03000593,
        64'h460943dc_fd843783,
        64'hdfc52781_8b89fe04,
        64'h2783a83d_fef42623,
        64'h4785c91f_f0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hc3852781_8ff967a1,
        64'hfe042703_fef42023,
        64'h87aac7ff_f0ef853e,
        64'h03000593_43dcfd84,
        64'h3783a8bd_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hc85fe0ef_fd843503,
        64'h30078593_67ad4601,
        64'h86be2781_fe645783,
        64'h7010d073_70105073,
        64'h0ff0000f_c2e19423,
        64'h4745ebcf_f0effd84,
        64'h350385be_fd043603,
        64'h2781fe64_5783d1df,
        64'hf0ef853e_4591863a,
        64'hfe445703_43dcfd84,
        64'h3783fef4_12238ff9,
        64'h17fd6785_fe445703,
        64'hfef41223_47a1fef4,
        64'h13234785_a201fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aad07f_e0effd84,
        64'h35037007_8593678d,
        64'h863e4681_4bbcfd84,
        64'h3783fce7_dfe3479d,
        64'h0007871b_fe842783,
        64'hfef42423_2785fe84,
        64'h27830007_802397ba,
        64'hfd043703_fe842783,
        64'haaa14785_c2e1a223,
        64'h4705ae6f_d0ef9365,
        64'h05130000_251792e5,
        64'h85930000_25970ba0,
        64'h0613a835_fe042423,
        64'hc201a223_a2514785,
        64'hc2e1a223_4705b12f,
        64'hd0ef9625_05130000,
        64'h251795a5_85930000,
        64'h25970b90_0613a015,
        64'h02f71963_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_c201a223,
        64'hcf91fd84_3783fcb4,
        64'h3823fca4_3c231800,
        64'hf022f406_71798082,
        64'h61457402_70a2853e,
        64'hfec42783_fe042623,
        64'he2fff0ef_85364591,
        64'h863e93c1_17c28ff9,
        64'h17fd6785_fd645703,
        64'h43d4fd84_3783fef4,
        64'h26232781_87aada9f,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfd84,
        64'h3783a081_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'he25fe0ef_fd843503,
        64'h6585863e_46812781,
        64'hfd645783_a0adfef4,
        64'h26234785_a89d4785,
        64'hc2e1a223_4705be2f,
        64'hd0efa325_05130000,
        64'h2517a2a5_85930000,
        64'h259707f0_0613a015,
        64'hc79d2781_3037f793,
        64'hfe842783_fef42423,
        64'h87aae25f_f0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'hc201a223_a0d94785,
        64'hc2e1a223_4705c32f,
        64'hd0efa825_05130000,
        64'h2517a7a5_85930000,
        64'h259707e0_0613a015,
        64'h04f71b63_11178793,
        64'h111117b7_873e53dc,
        64'hfd843783_c201a223,
        64'hcf91fd84_3783fcf4,
        64'h1b2387ae_fca43c23,
        64'h1800f022_f4067179,
        64'h80826105_644260e2,
        64'h0001eb7f_f0ef853e,
        64'h85bafea4_47039381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef40523_87bafef4,
        64'h05a387b6_fef42623,
        64'h873286ae_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e2853e,
        64'h87aaea9f_f0ef853e,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_05a387ba,
        64'hfef42623_872e87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h0001f63f_f0ef853e,
        64'h85bafe84_57039381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef41423_87bafef4,
        64'h05a387b6_fef42623,
        64'h873286ae_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e2853e,
        64'h87aaf47f_f0ef853e,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_05a387ba,
        64'hfef42623_872e87aa,
        64'h1000e822_ec061101,
        64'h80826145_74220001,
        64'h00e79023_fd645703,
        64'hfe843783_fef43423,
        64'hfd843783_fcf41b23,
        64'h87aefca4_3c231800,
        64'hf4227179_80826145,
        64'h74220001_00e78023,
        64'hfd744703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf40ba3_87aefca4,
        64'h3c231800_f4227179,
        64'h80826105_6462853e,
        64'h2781439c_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61056462,
        64'h853e93c1_17c20007,
        64'hd783fe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826105_6462853e,
        64'h0ff7f793_0007c783,
        64'hfe843783_fea43423,
        64'h1000ec22_11018082,
        64'h61616406_60a6853e,
        64'hfec42783_fe042623,
        64'hd3f8fb84_37830007,
        64'h871b0097_d79bfd84,
        64'h2783fcf4_2c2302f7,
        64'h07bbfe04_2783fd84,
        64'h2703fcf4_2c2302f7,
        64'h07bbfdc4_27032781,
        64'h2785fd84_2783fcf4,
        64'h2c238fd9_fd842783,
        64'h0007871b_8ff9c007,
        64'h87936785_873e2781,
        64'h00a7979b_fd042783,
        64'hfcf42c23_0167d79b,
        64'hfcc42783_fcf42e23,
        64'h278100f7_17bb4705,
        64'h27812789_27818b9d,
        64'h27810077_d79bfcc4,
        64'h2783fef4_20232781,
        64'h00f717bb_47052781,
        64'h8bbd2781_0087d79b,
        64'hfd042783_02e78aa3,
        64'hfb843783_0ff7f713,
        64'h8bbd0ff7_f7932781,
        64'h0127d79b_fd442783,
        64'hfcf42a23_278187aa,
        64'ha11fd0ef_853e9381,
        64'h17822781_27f143dc,
        64'hfb843783_fcf42823,
        64'h278187aa_a2dfd0ef,
        64'h853e9381_17822781,
        64'h27e143dc_fb843783,
        64'hfcf42623_278187aa,
        64'ha49fd0ef_853e9381,
        64'h17822781_27d143dc,
        64'hfb843783_fcf42423,
        64'h278187aa_a65fd0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fb843783,
        64'ha23dfef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa9e2f,
        64'hf0effb84_35039007,
        64'h85936785_863e4681,
        64'h4bbcfb84_3783aab1,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_a10ff0ef,
        64'hfb843503_30000593,
        64'h863e4681_4bbcfb84,
        64'h3783cbb8_12340737,
        64'hfb843783_c7f8fb84,
        64'h37830007_871b87aa,
        64'hb85fd0ef_853e45f1,
        64'h43dcfb84_3783c7b8,
        64'hfb843783_0007871b,
        64'h87aab9ff_d0ef853e,
        64'h45e143dc_fb843783,
        64'hc3f8fb84_37830007,
        64'h871b87aa_bb9fd0ef,
        64'h853e45d1_43dcfb84,
        64'h3783c3b8_fb843783,
        64'h0007871b_87aabd3f,
        64'hd0ef853e_45c143dc,
        64'hfb843783_aaedfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaaaef_f0effb84,
        64'h35032000_05934601,
        64'h4681db98_4705fb84,
        64'h3783c789_27818ff9,
        64'h400007b7_fe842703,
        64'hfa07dde3_fe842783,
        64'hfef42423_87aab8ff,
        64'hd0ef853e_93811782,
        64'h278127c1_43dcfb84,
        64'h3783aca1_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'hb0cff0ef_fb843503,
        64'h10000593_40ff8637,
        64'h4681a091_fe042423,
        64'ha459fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aab3af,
        64'hf0effb84_35034581,
        64'h46014681_a46dfef4,
        64'h26234785_e7892781,
        64'h8ff967c1_fe442703,
        64'hfef42223_87aac0ff,
        64'hd0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfb843783_cb8d47dc,
        64'hfb843783_02f70e63,
        64'h400007b7_873e2781,
        64'h8ff9c000_07b7873e,
        64'h579cfb84_3783a601,
        64'h4785c2e1_a2234705,
        64'h93dfd0ef_f6c50513,
        64'h00002517_f6c58593,
        64'h00002597_68900613,
        64'ha01504f7_11634789,
        64'h873e0367_c783fb84,
        64'h3783c201_a223ae25,
        64'h4785c2e1_a2234705,
        64'h975fd0ef_fa450513,
        64'h00002517_fa458593,
        64'h00002597_68800613,
        64'ha01502f7_1f631117,
        64'h87931111_17b7873e,
        64'h53dcfb84_3783c201,
        64'ha223cf91_fb843783,
        64'hfaa43c23_0880e0a2,
        64'he486715d_80826121,
        64'h744270e2_00017010,
        64'hd0737010_50730ff0,
        64'h000fd55f_d0ef853a,
        64'h85be2781_08078793,
        64'hfd843783_93010207,
        64'h97132781_0587879b,
        64'h43dcfd84_378300e7,
        64'h912397b6_078e07c1,
        64'h93810206_1793fd84,
        64'h36839341_03079713,
        64'h02f707bb_0006861b,
        64'h36fdfec4_268393c1,
        64'h17c2fe44_27839341,
        64'h03079713_fd442783,
        64'h00e79023_02300713,
        64'h97ba078e_07c19381,
        64'h1782fd84_37032781,
        64'h37fdfec4_2783c3d8,
        64'h97b6078e_07c19381,
        64'h02061793_fd843683,
        64'h0007871b_9fb90006,
        64'h861b36fd_fec42683,
        64'h27810107_979bfe84,
        64'h27830007_871bfc84,
        64'h3783f8e7_ebe32781,
        64'hfe842783_0007871b,
        64'h37fdfec4_2783fef4,
        64'h24232785_fe842783,
        64'h00079123_97ba078e,
        64'h07c1fe84_6783fd84,
        64'h370300e7_90230210,
        64'h071397ba_078e07c1,
        64'hfe846783_fd843703,
        64'hc3d897b6_078e07c1,
        64'hfe846783_fd843683,
        64'h0007871b_9fb92781,
        64'h0107979b_fe842783,
        64'h0007871b_fc843783,
        64'ha8b1fe04_2423fef4,
        64'h26232785_fec42783,
        64'hc7912781_8ff917fd,
        64'h67c1873e_278102f7,
        64'h07bbfe44_2783fd44,
        64'h2703fef4_26230107,
        64'hd79b2781_02f707bb,
        64'hfe442783_fd442703,
        64'ha835fef4_26234785,
        64'h00f77663_67c1873e,
        64'h278102f7_07bbfe44,
        64'h2783fd44_2703fef4,
        64'h22238ff9_17fd6785,
        64'hfe442703_fef42223,
        64'h87aaf0ff_d0ef853e,
        64'h459143dc_fd843783,
        64'hfe042223_fe042423,
        64'hfe042623_fcf42a23,
        64'hfcc43423_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_61457402,
        64'h70a2853e_fec42783,
        64'h0001a011_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'he1cff0ef_fd843503,
        64'h70000593_863e4681,
        64'h4bbcfd84_3783fe04,
        64'h2623fca4_3c231800,
        64'hf022f406_71798082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hfd7fd0ef_853e0300,
        64'h05934609_43dcfd84,
        64'h3783dfc5_27818b89,
        64'hfe442783_a00dfef4,
        64'h26234785_ffbfd0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_fe9fd0ef,
        64'h853e0300_059343dc,
        64'hfd843783_a08dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aaec6f_f0effd84,
        64'h35039007_85936789,
        64'h863e86ba_fd442783,
        64'hfd042703_c2e19423,
        64'h02700713_a869fef4,
        64'h26234785_c3a92781,
        64'hfec42783_fef42623,
        64'h87aaefef_f0effd84,
        64'h35038007_85936789,
        64'h863e86ba_fd442783,
        64'hfd042703_c2e19423,
        64'h470d02f7_1d634785,
        64'h0007871b_fd042783,
        64'h7010d073_70105073,
        64'h0ff0000f_146000ef,
        64'hfd843503_85befc84,
        64'h3603fd04_2783a8f5,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_081000ef,
        64'hfd843503_20000593,
        64'h02f70363_20000793,
        64'h873e2781_87aa826f,
        64'he0ef853e_93811782,
        64'h27812791_43dcfd84,
        64'h3783a281_fef42623,
        64'h4785e789_27818ff9,
        64'h67c1fe84_2703fef4,
        64'h242387aa_854fe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783cb8d_47dcfd84,
        64'h378302f7_0e634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfd843783_00f71f63,
        64'h4789873e_0367c783,
        64'hfd843783_fcf42823,
        64'h87bafcf4_2a23fcd4,
        64'h34238732_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_61217442,
        64'h70e2853e_fec42783,
        64'hfe042623_fef42623,
        64'h278187aa_8d4fe0ef,
        64'h853e9381_17822781,
        64'h27c143dc_fd843783,
        64'h9befe0ef_853e0300,
        64'h05934609_43dcfd84,
        64'h3783dfc5_27818b89,
        64'hfe442783_a83dfef4,
        64'h26234785_9e2fe0ef,
        64'h853a0320_05933ff7,
        64'h861367bd_43d8fd84,
        64'h3783c385_27818ff9,
        64'h67a1fe44_2703fef4,
        64'h222387aa_9d0fe0ef,
        64'h853e0300_059343dc,
        64'hfd843783_a8bdfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa8aff_f0effd84,
        64'h35032007_85936785,
        64'h863e86ba_fd442783,
        64'hfd042703_c2e19423,
        64'h03700713_a85dfef4,
        64'h26234785_c3a92781,
        64'hfec42783_fef42623,
        64'h87aa8e7f_f0effd84,
        64'h35031007_85936785,
        64'h863e86ba_fd442783,
        64'hfd042703_c2e19423,
        64'h474d02f7_1d634785,
        64'h0007871b_fd042783,
        64'h7010d073_70105073,
        64'h0ff0000f_32e000ef,
        64'hfd843503_85befc84,
        64'h3603fd04_2783aa21,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_269000ef,
        64'hfd843503_20000593,
        64'h02f70363_20000793,
        64'h873e2781_87aaa0ef,
        64'he0ef853e_93811782,
        64'h27812791_43dcfd84,
        64'h3783aab1_fef42623,
        64'h4785e789_27818ff9,
        64'h67c1fe84_2703fef4,
        64'h242387aa_a3cfe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783cb8d_47dcfd84,
        64'h378302f7_0e634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfd843783_00f71f63,
        64'h4789873e_0367c783,
        64'hfd843783_fcf42823,
        64'h87bafcf4_2a23fcd4,
        64'h34238732_87aefca4,
        64'h3c230080_f822fc06,
        64'h71398082_61457422,
        64'h853efec4_27830001,
        64'ha0110001_a0210001,
        64'ha031fef4_26238fd9,
        64'hfd442783_fec42703,
        64'ha831fef4_262301a7,
        64'he793fec4_2783a02d,
        64'hfef42623_03a7e793,
        64'hfec42783_a825fef4,
        64'h262301a7_e793fec4,
        64'h2783a099_fef42623,
        64'h0027e793_fec42783,
        64'ha891fef4_262303a7,
        64'he793fec4_2783a08d,
        64'hfef42623_03a7e793,
        64'hfec42783_a885fef4,
        64'h262301a7_e793fec4,
        64'h2783a8bd_fef42623,
        64'h0097e793_fec42783,
        64'ha071fef4_262303a7,
        64'he793fec4_2783a869,
        64'hfef42623_01a7e793,
        64'hfec42783_00f71963,
        64'h4785873e_0347c783,
        64'hfd843783_a865fef4,
        64'h262301a7_e793fec4,
        64'h2783a0d9_fef42623,
        64'h01a7e793_fec42783,
        64'ha8d1fef4_262301b7,
        64'he793fec4_2783a0cd,
        64'hfef42623_03a7e793,
        64'hfec42783_00f71963,
        64'h4785873e_0347c783,
        64'hfd843783_a201fef4,
        64'h262301b7_e793fec4,
        64'h2783a239_fef42623,
        64'h01b7e793_fec42783,
        64'haa31fef4_26230097,
        64'he793fec4_2783a22d,
        64'hfef42623_0027e793,
        64'hfec42783_aa390ef7,
        64'h05639007_879367ad,
        64'h0007871b_10e68a63,
        64'h30070713_672d0007,
        64'h869b10e6_8a63a007,
        64'h0713672d_0007869b,
        64'ha2a916f7_0363a007,
        64'h87936791_0007871b,
        64'h0ee68d63_d0070713,
        64'h67250007_869b0ae6,
        64'h89636007_07136721,
        64'h0007869b_02d76863,
        64'h70070713_67250007,
        64'h869b14e6_80637007,
        64'h07136725_0007869b,
        64'haa4914f7_08638007,
        64'h87936789_0007871b,
        64'h18e68b63_40070713,
        64'h670d0007_869b16e6,
        64'h86639007_07136709,
        64'h0007869b_aa7d16f7,
        64'h07632007_87936785,
        64'h0007871b_16e68e63,
        64'h50070713_67050007,
        64'h869b18e6_85633007,
        64'h07136705_0007869b,
        64'h02d76863_70070713,
        64'h67050007_869b1ae6,
        64'h8a637007_07136705,
        64'h0007869b_06d76c63,
        64'h70070713_670d0007,
        64'h869b20e6_84637007,
        64'h0713670d_0007869b,
        64'ha40d1cf7_0263b007,
        64'h87936785_0007871b,
        64'h1ce68963_67050007,
        64'h869b1ce6_8e63c007,
        64'h07136705_0007869b,
        64'ha4a91af7_02637000,
        64'h07930007_871b1ee6,
        64'h85639007_07136705,
        64'h0007869b_1c070663,
        64'h27018007_871b02d7,
        64'h6563a007_07136705,
        64'h0007869b_20e68f63,
        64'ha0070713_67050007,
        64'h869ba471_18f70863,
        64'h30000793_0007871b,
        64'h1ae68563_50000713,
        64'h0007869b_2ae68e63,
        64'h40000713_0007869b,
        64'hac4d18f7_0d631000,
        64'h07930007_871b2c07,
        64'h09630007_871b00d7,
        64'h6d632000_07130007,
        64'h869b1ce6_84632000,
        64'h07130007_869b04d7,
        64'h6c636000_07130007,
        64'h869b20e6_85636000,
        64'h07130007_869b0cd7,
        64'h6d631007_07136705,
        64'h0007869b_2ae68a63,
        64'h10070713_67050007,
        64'h869bfd44_2783fef4,
        64'h2623fd44_2783fcf4,
        64'h2a2387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61217442_70e2853e,
        64'hfec42783_fe042623,
        64'hedefe0ef_853e0300,
        64'h05934605_43dcfd84,
        64'h3783d3a9_27818b85,
        64'hfe042783_a00defcf,
        64'he0ef853a_03200593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_fef42623,
        64'h4789e781_27819bf9,
        64'hfec42783_fef42623,
        64'h87aaeeef_e0ef853e,
        64'h03200593_43dcfd84,
        64'h3783c3a1_27818ff9,
        64'h67a1fe04_2703a899,
        64'hf46fe0ef_853e0300,
        64'h05930200_061343dc,
        64'hfd843783_cf812781,
        64'h0207f793_278187aa,
        64'hf2cfe0ef_853e0300,
        64'h059343dc_fd843783,
        64'h02f71b63_30078793,
        64'h67850007_871bfd44,
        64'h278300f7_0b635007,
        64'h87936785_0007871b,
        64'hfd442783_fef42023,
        64'h87aaf66f_e0ef853e,
        64'h03000593_43dcfd84,
        64'h3783f4cf_e0ef853a,
        64'h85be2781_8fd52781,
        64'hc281d783_0007869b,
        64'h0107979b_fe442783,
        64'h93010207_97132781,
        64'h27b143dc_fd843783,
        64'ha219fef4_26234785,
        64'hc7892781_0207f793,
        64'hfe442783_cb992781,
        64'h8b89fe84_2783fef4,
        64'h242387aa_f2cfe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h378302f7_0f633007,
        64'h87936785_0007871b,
        64'hfd442783_04f70863,
        64'h50078793_67850007,
        64'h871bfd44_2783fef4,
        64'h22238ff9_17fd6791,
        64'hfe442703_fef42223,
        64'h87aa1880_00effd84,
        64'h350385be_fd442783,
        64'h85ffe0ef_853a0320,
        64'h05933ff7_861367bd,
        64'h43d8fd84_3783875f,
        64'he0ef853a_03000593,
        64'hfff78613_67c143d8,
        64'hfd843783_827fe0ef,
        64'h853e85ba_fd042703,
        64'h93811782_278127a1,
        64'h43dcfd84_3783925f,
        64'he0ef853e_02e00593,
        64'h463943dc_fd843783,
        64'h8b7fe0ef_853e4599,
        64'h863a9341_1742fcc4,
        64'h270343dc_fd843783,
        64'haaddfef4_26234785,
        64'ha4094785_c2e1a223,
        64'h4705cf6f_e0efb265,
        64'h05130000_3517b265,
        64'h85930000_359744c0,
        64'h0613a015_c79d2781,
        64'h8b85fe84_2783fef4,
        64'h242387aa_835fe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783c201_a223ac81,
        64'h4785c2e1_a2234705,
        64'hd44fe0ef_b7450513,
        64'h00003517_b7458593,
        64'h00003597_44b00613,
        64'ha01504f7_1a631117,
        64'h87931111_17b7873e,
        64'h53dcfd84_3783c201,
        64'ha223cf91_fd843783,
        64'hfcf42623_87bafcf4,
        64'h282387b2_fcf42a23,
        64'h873687ae_fca43c23,
        64'h0080f822_fc067139,
        64'h80826145_740270a2,
        64'h853efec4_27830001,
        64'hfcf719e3_01f007b7,
        64'h873e2781_8ff901f0,
        64'h07b7fe84_2703fef4,
        64'h242387aa_8ddfe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783a839_fef42423,
        64'h87aa8fbf_e0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fd843783,
        64'h80ffe0ef_3e800513,
        64'h9effe0ef_853a02c0,
        64'h0593863e_93c117c2,
        64'h0047e793_93c117c2,
        64'hfe442783_43d8fd84,
        64'h3783fef4_222387aa,
        64'h9ddfe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'hd3ed2781_8b89fe44,
        64'h2783fef4_222387aa,
        64'h9fdfe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'ha821fef4_222387aa,
        64'ha15fe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'ha5ffe0ef_853a02c0,
        64'h0593863e_93c117c2,
        64'h0017e793_93c117c2,
        64'hfe442783_43d8fd84,
        64'h3783fef4_222387aa,
        64'ha4dfe0ef_853e02c0,
        64'h059343dc_fd843783,
        64'ha211fef4_26234785,
        64'he7892781_8ba12781,
        64'hfe245783_fef41123,
        64'h87aaa77f_e0ef853e,
        64'h03e00593_43dcfd84,
        64'h37838e9f_e0ef3887,
        64'h85136785_acbfe0ef,
        64'h853e03e0_0593863a,
        64'hfe245703_43dcfd84,
        64'h3783fef4_11230087,
        64'he793fe24_5783fef4,
        64'h112387aa_ab9fe0ef,
        64'h853e03e0_059343dc,
        64'hfd843783_b03fe0ef,
        64'h853e02c0_0593863a,
        64'hfe245703_43dcfd84,
        64'h3783fef4_11239be9,
        64'hfe245783_fef41123,
        64'h87aaaeff_e0ef853e,
        64'h02c00593_43dcfd84,
        64'h3783ffe1_27818ff9,
        64'h01f007b7_fe842703,
        64'hfef42423_87aaa77f,
        64'he0ef853e_93811782,
        64'h27810247_879b43dc,
        64'hfd843783_a839fef4,
        64'h242387aa_a95fe0ef,
        64'h853e9381_17822781,
        64'h0247879b_43dcfd84,
        64'h3783fef4_26234785,
        64'hc7812781_fec42783,
        64'hfef42623_87aa2120,
        64'h00effd84_3503b007,
        64'h85936785_46014681,
        64'hfca43c23_1800f022,
        64'hf4067179_80826145,
        64'h740270a2_853efec4,
        64'h2783fe04_2623f3e5,
        64'h27818b89_2781feb4,
        64'h4783fef4_05a387aa,
        64'hc1dfe0ef_853e02f0,
        64'h059343dc_fd843783,
        64'ha821fef4_05a387aa,
        64'hc35fe0ef_853e02f0,
        64'h059343dc_fd843783,
        64'hc7ffe0ef_853e02f0,
        64'h05934609_43dcfd84,
        64'h3783c11f_e0ef853a,
        64'h03200593_3ff78613,
        64'h67bd43d8_fd843783,
        64'hc27fe0ef_853a0300,
        64'h0593fff7_861367c1,
        64'h43d8fd84_378302e7,
        64'h8a234709_fd843783,
        64'ha03102e7_8a234705,
        64'hfd843783_c7992781,
        64'hfec42783_fef42623,
        64'h87aa2de0_00effd84,
        64'h35031000_059340ff,
        64'h86374681_a855fef4,
        64'h26234785_a0c14785,
        64'hc2e1a223_470589bf,
        64'he0efeca5_05130000,
        64'h3517eca5_85930000,
        64'h35973ac0_0613a015,
        64'hc79d2781_fec42783,
        64'hfef42623_87aa32a0,
        64'h00effd84_35034581,
        64'h46014681_ae3fe0ef,
        64'h71078513_6789c201,
        64'ha223a239_4785c2e1,
        64'ha2234705_8e9fe0ef,
        64'hf1850513_00003517,
        64'hf1858593_00003597,
        64'h3ab00613_a01504f7,
        64'h1a631117_87931111,
        64'h17b7873e_53dcfd84,
        64'h3783c201_a223cf91,
        64'hfd843783_fca43c23,
        64'h1800f022_f4067179,
        64'h8082614d_64ea740a,
        64'h70aa853e_fdc42783,
        64'h0001a011_0001a021,
        64'h0001a031_fcf42e23,
        64'h4785cb89_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h4e4010ef_f5843503,
        64'h20000593_02f71763,
        64'h4785873e_0347c783,
        64'hf5843783_00f71a63,
        64'h4791873e_57fcf584,
        64'h37830001_a0b9fcf4,
        64'h2e234785_c7912781,
        64'hfdc42783_fcf42e23,
        64'h87aa71e0_20eff584,
        64'h350385be_fd442783,
        64'hfcf42a23_1007879b,
        64'h03a207b7_eb950a27,
        64'hc78307a7_87931ffe,
        64'hd797a071_fcf42e23,
        64'h4785c789_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h065010ef_f5843503,
        64'h02f71163_4791873e,
        64'h57fcf584_3783a865,
        64'hfcf42e23_478500f7,
        64'h06634785_873e0b97,
        64'hc7830c27_87931ffe,
        64'hd79704f7_16634791,
        64'h873e57fc_f5843783,
        64'h00f70963_4795873e,
        64'h57fcf584_3783a8c5,
        64'hfcf42e23_478500f7,
        64'h06634789_873e0b97,
        64'hc7830fa7_87931ffe,
        64'hd79702f7_1063479d,
        64'h873e57fc_f5843783,
        64'haa29fcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa6340,
        64'h20eff584_350312e5,
        64'h85931ffe_d597a281,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_607010ef,
        64'hf5843503_0cf70b63,
        64'h4799873e_57fcf584,
        64'h3783d7f8_4719f584,
        64'h3783a029_d7f84715,
        64'hf5843783_00e7f763,
        64'h4785873e_0377c783,
        64'hf5843783_cf912781,
        64'h8b892781_0c47c783,
        64'h19078793_1ffed797,
        64'ha825d7f8_4711f584,
        64'h378300e7_f7634785,
        64'h873e0377_c783f584,
        64'h3783cf91_27818bb1,
        64'h27810c47_c7831be7,
        64'h87931ffe_d797a09d,
        64'hd7f8471d_f5843783,
        64'h00e7f763_4785873e,
        64'h0377c783_f5843783,
        64'hcf912781_0307f793,
        64'h27810c47_c7831ee7,
        64'h87931ffe_d797d3f8,
        64'hf5843783_0007871b,
        64'h8fd92781_0d47c783,
        64'h20878793_1ffed797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h8fd92781_0087979b,
        64'h27810d57_c78322e7,
        64'h87931ffe_d79753f8,
        64'hf5843783_d3f8f584,
        64'h37830007_871b8fd9,
        64'h27810107_979b2781,
        64'h0d67c783_25478793,
        64'h1ffed797_53f8f584,
        64'h3783d3f8_f5843783,
        64'h0007871b_0187979b,
        64'h27810d77_c7832767,
        64'h87931ffe_d797a461,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_7a2020ef,
        64'hf5843503_29c58593,
        64'h1ffed597_a47dfcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa2870_10eff584,
        64'h350328f7_12634795,
        64'h873e0347_c783f584,
        64'h3783acf1_fcf42e23,
        64'h478528f7_0d634785,
        64'h873e0b97_c7832e67,
        64'h87931ffe_d797ace5,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_013020ef,
        64'hf5843503_30c58593,
        64'h1ffed597_ae39fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa7e50_10eff584,
        64'h3503d7f8_4715f584,
        64'h37832ee7_fd634785,
        64'h873e0377_c783f584,
        64'h37833007_85632781,
        64'h8b892781_0c47c783,
        64'h35878793_1ffed797,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810d47,
        64'hc7833727_87931ffe,
        64'hd79753f8_f5843783,
        64'hd3f8f584_37830007,
        64'h871b8fd9_27810087,
        64'h979b2781_0d57c783,
        64'h39878793_1ffed797,
        64'h53f8f584_3783d3f8,
        64'hf5843783_0007871b,
        64'h8fd92781_0107979b,
        64'h27810d67_c7833be7,
        64'h87931ffe_d79753f8,
        64'hf5843783_d3f8f584,
        64'h37830007_871b0187,
        64'h979b2781_0d77c783,
        64'h3e078793_1ffed797,
        64'haecdfcf4_2e234785,
        64'hc7892781_fdc42783,
        64'hfcf42e23_87aa10d0,
        64'h20eff584_35034065,
        64'h85931ffe_d597a921,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_3f1010ef,
        64'hf5843503_14f71f63,
        64'h4785873e_0367c783,
        64'hf5843783_16e7f763,
        64'h478d873e_0357c783,
        64'hf5843783_16f71f63,
        64'h4789873e_0347c783,
        64'hf5843783_a19dfcf4,
        64'h2e234785_42078363,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_12e020ef,
        64'hf5843503_d7f84715,
        64'hf5843783_44e7f363,
        64'h4785873e_0377c783,
        64'hf5843783_44078b63,
        64'h27818b89_2781f9d4,
        64'h47834607_82630004,
        64'hc78302e7_8e234705,
        64'hf5843783_80aff0ef,
        64'h3e800513_9eaff0ef,
        64'h853a02c0_0593863e,
        64'h93c117c2_0047e793,
        64'hfda45783_43d8f584,
        64'h3783fcf4_1d2387aa,
        64'h9d4ff0ef_853e02c0,
        64'h059343dc_f5843783,
        64'hd3e52781_8b892781,
        64'hfda45783_fcf41d23,
        64'h87aa9f6f_f0ef853e,
        64'h02c00593_43dcf584,
        64'h3783a821_fcf41d23,
        64'h87aaa0ef_f0ef853e,
        64'h02c00593_43dcf584,
        64'h3783a58f_f0ef853a,
        64'h02c00593_863e93c1,
        64'h17c20017_e793fda4,
        64'h578343d8_f5843783,
        64'hfcf41d23_87aaa42f,
        64'hf0ef853e_02c00593,
        64'h43dcf584_3783a3a5,
        64'hfcf42e23_4785e789,
        64'h27818ba1_2781fd24,
        64'h5783fcf4_192387aa,
        64'ha6cff0ef_853e03e0,
        64'h059343dc_f5843783,
        64'h8deff0ef_38878513,
        64'h6785ac0f_f0ef853e,
        64'h03e00593_863afd24,
        64'h570343dc_f5843783,
        64'hfcf41923_0087e793,
        64'hfd245783_fcf41923,
        64'h87aaaaef_f0ef853e,
        64'h03e00593_43dcf584,
        64'h3783af8f_f0ef853e,
        64'h02c00593_863afd24,
        64'h570343dc_f5843783,
        64'hfcf41923_9be9fd24,
        64'h5783fcf4_192387aa,
        64'hae4ff0ef_853e02c0,
        64'h059343dc_f5843783,
        64'h14079d63_03c7c783,
        64'hf5843783_16f71363,
        64'h47a1873e_4bdcf584,
        64'h378316e7_fa63478d,
        64'h873ef9d4_47831807,
        64'hd0634187_d79b0187,
        64'h979b0024_c7836207,
        64'h9e632781_fdc42783,
        64'hfcf42e23_87aa1460,
        64'h20eff584_350385be,
        64'hf9040793_adb9fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa6370_10eff584,
        64'h3503c385_27818b91,
        64'h27810014_c783a561,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_483010ef,
        64'hf5843503_85a6a565,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_2e5020ef,
        64'hf5843503_26f71263,
        64'h4785873e_0347c783,
        64'hf5843783_add9fcf4,
        64'h2e234785_c7892781,
        64'hfdc42783_fcf42e23,
        64'h87aa4500_10eff584,
        64'h3503add5_fcf42e23,
        64'h4785adf5_fcf42e23,
        64'h4785cb89_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h017020ef_f5843503,
        64'h85be5f9c_f5843783,
        64'hdf98a807_071b018c,
        64'hc737f584_3783af05,
        64'hfcf42e23_4785c789,
        64'h2781fdc4_2783fcf4,
        64'h2e2387aa_6cc010ef,
        64'hf5843503_04f71b63,
        64'h4795873e_0347c783,
        64'hf5843783_00f70a63,
        64'h4789873e_0347c783,
        64'hf5843783_a7bdfcf4,
        64'h2e234785_c3d12781,
        64'hfdc42783_fcf42e23,
        64'h87aa0890_20eff584,
        64'h350385be_5f9cf584,
        64'h3783df98_8407071b,
        64'h017d8737_f5843783,
        64'ha801df98_ac07071b,
        64'h0121f737_f5843783,
        64'h00f71a63_4789873e,
        64'h0367c783_f5843783,
        64'h7c40006f_fcf42e23,
        64'h4785c791_2781fdc4,
        64'h2783fcf4_2e2387aa,
        64'h935ff0ef_f5843503,
        64'h06f71c63_4785873e,
        64'h0347c783_f5843783,
        64'h7f40006f_fcf42e23,
        64'h478500f7_07634795,
        64'h873e0347_c783f584,
        64'h378300f7_0f634789,
        64'h873e0347_c783f584,
        64'h378302f7_07634785,
        64'h873e0347_c783f584,
        64'h378302f7_02e34785,
        64'h0007871b_fdc42783,
        64'hfcf42e23_87aa0530,
        64'h00eff584_3503a839,
        64'h02e78a23_4715f584,
        64'h378300f7_18634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hf5843783_0750006f,
        64'h4785c2e1_a2234705,
        64'h9b4ff0ef_7e450513,
        64'h00003517_7e458593,
        64'h00003597_24000613,
        64'ha01d04f7_18634789,
        64'h873e0367_c783f584,
        64'h3783df98_a807071b,
        64'h00062737_f5843783,
        64'h02078e23_f5843783,
        64'h02e78a23_4705f584,
        64'h378302e7_8ba34705,
        64'hf5843783_c201a223,
        64'h0d90006f_4785c2e1,
        64'ha2234705_a18ff0ef,
        64'h84850513_00004517,
        64'h84858593_00004597,
        64'h23f00613_a01d06f7,
        64'h15631117_87931111,
        64'h17b7873e_53dcf584,
        64'h3783c201_a223cf91,
        64'hf5843783_fc043423,
        64'hfc043023_fa043c23,
        64'hfa043823_fa043423,
        64'hfa043023_f8043c23,
        64'hf8043823_0004b023,
        64'h00579493_839507fd,
        64'hf8078793_fe040793,
        64'hf4a43c23_1900ed26,
        64'hf122f506_71718082,
        64'h61616406_60a6853e,
        64'hfec42783_fe042623,
        64'hd3f8fb84_37830007,
        64'h871b00a7_979b2781,
        64'h27852781_8ff917fd,
        64'h004007b7_873e2781,
        64'h0087d79b_fc442783,
        64'h02f71663_4785873e,
        64'h27818b8d_27810167,
        64'hd79bfcc4_2783a081,
        64'hd3f8fb84_37830007,
        64'h871b0097_d79bfd04,
        64'h2783fcf4_282302f7,
        64'h07bbfd84_2783fd04,
        64'h2703fcf4_282302f7,
        64'h07bbfd44_27032781,
        64'h2785fd04_2783fcf4,
        64'h28238fd9_fd042783,
        64'h0007871b_8ff9c007,
        64'h87936785_873e2781,
        64'h00a7979b_fc842783,
        64'hfcf42823_0167d79b,
        64'hfc442783_fcf42a23,
        64'h278100f7_17bb4705,
        64'h27812789_27818b9d,
        64'h27810077_d79bfc44,
        64'h2783fcf4_2c232781,
        64'h00f717bb_47052781,
        64'h8bbd2781_0087d79b,
        64'hfc842783_e3c52781,
        64'h8b8d2781_0167d79b,
        64'hfcc42783_fcf42623,
        64'h278187aa_eacff0ef,
        64'h853e9381_17822781,
        64'h27f143dc_fb843783,
        64'hfcf42423_278187aa,
        64'hec8ff0ef_853e9381,
        64'h17822781_27e143dc,
        64'hfb843783_fcf42223,
        64'h278187aa_ee4ff0ef,
        64'h853e9381_17822781,
        64'h27d143dc_fb843783,
        64'hfcf42023_278187aa,
        64'hf00ff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_a28dfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa67f0_00effb84,
        64'h35039007_85936785,
        64'h863e4681_4bbcfb84,
        64'h3783d7d5_4bbcfb84,
        64'h3783cbb8_fb843783,
        64'h0007871b_8ff977c1,
        64'h873e2781_87aaf5ef,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfb84,
        64'h3783a2c1_fef42623,
        64'h4785c789_2781fec4,
        64'h2783fef4_262387aa,
        64'h6dd000ef_fb843503,
        64'h30000593_46014681,
        64'hc7f8fb84_37830007,
        64'h871b87aa_841ff0ef,
        64'h853e45f1_43dcfb84,
        64'h3783c7b8_fb843783,
        64'h0007871b_87aa85bf,
        64'hf0ef853e_45e143dc,
        64'hfb843783_c3f8fb84,
        64'h37830007_871b87aa,
        64'h875ff0ef_853e45d1,
        64'h43dcfb84_3783c3b8,
        64'hfb843783_0007871b,
        64'h87aa88ff_f0ef853e,
        64'h45c143dc_fb843783,
        64'ha4b9fef4_26234785,
        64'hc7892781_fec42783,
        64'hfef42623_87aa76b0,
        64'h00effb84_35032000,
        64'h05934601_4681ac95,
        64'hfef42623_4785c789,
        64'h2781fec4_2783fef4,
        64'h262387aa_565000ef,
        64'hfb843503_02e78e23,
        64'h4705fb84_3783c78d,
        64'h27818ff9_010007b7,
        64'hfe842703_db984705,
        64'hfb843783_c7892781,
        64'h8ff94000_07b7fe84,
        64'h2703f407_dde3fe84,
        64'h2783fef4_242387aa,
        64'h881ff0ef_853e9381,
        64'h17822781_27c143dc,
        64'hfb843783_a4cdfef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa7ff0_00effb84,
        64'h35039007_859367ad,
        64'h863e4681_fe442783,
        64'hfef42223_8fd90100,
        64'h07b7fe44_270300f7,
        64'h196347a1_873e4bdc,
        64'hfb843783_02f71063,
        64'h4789873e_0367c783,
        64'hfb843783_fef42223,
        64'h40ff87b7_a689fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa05e0_10effb84,
        64'h35037007_8593678d,
        64'h46014681_a055fe04,
        64'h242302e7_8aa34709,
        64'hfb843783_a03102e7,
        64'h8aa34705_fb843783,
        64'h00f70863_1aa00793,
        64'h0007871b_fe842783,
        64'hfef42423_87aa94ff,
        64'hf0ef853e_93811782,
        64'h278127c1_43dcfb84,
        64'h3783f3e5_27818b89,
        64'h2781fe34_4783fef4,
        64'h01a387aa_a91ff0ef,
        64'h853e02f0_059343dc,
        64'hfb843783_a821fef4,
        64'h01a387aa_aa9ff0ef,
        64'h853e02f0_059343dc,
        64'hfb843783_af3ff0ef,
        64'h853e02f0_05934609,
        64'h43dcfb84_378304f7,
        64'h18634789_0007871b,
        64'hfec42783_a129fef4,
        64'h26234785_00f70663,
        64'h47890007_871bfec4,
        64'h2783cf81_2781fec4,
        64'h2783fef4_262387aa,
        64'h134010ef_fb843503,
        64'h80078593_67851aa0,
        64'h06134681_a189fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa15e0_10effb84,
        64'h35034581_46014681,
        64'ha19dfef4_26234785,
        64'he7892781_8ff967c1,
        64'hfdc42703_fcf42e23,
        64'h87aaa33f_f0ef853e,
        64'h93811782_27810247,
        64'h879b43dc_fb843783,
        64'hcb8d47dc_fb843783,
        64'h02f70e63_400007b7,
        64'h873e2781_8ff9c000,
        64'h07b7873e_579cfb84,
        64'h3783a975_4785c2e1,
        64'ha2234705_f60ff0ef,
        64'hd9050513_00004517,
        64'hd9058593_00004597,
        64'h16200613_a01504f7,
        64'h11634789_873e0367,
        64'hc783fb84_3783cbd8,
        64'h4711fb84_3783c201,
        64'ha223a9f5_4785c2e1,
        64'ha2234705_fa0ff0ef,
        64'hdd050513_00004517,
        64'hdd058593_00004597,
        64'h16100613_a01504f7,
        64'h13631117_87931111,
        64'h17b7873e_53dcfb84,
        64'h3783c201_a223cf91,
        64'hfb843783_faa43c23,
        64'h0880e0a2_e486715d,
        64'h80826121_744270e2,
        64'h853efec4_2783fe04,
        64'h2623be1f_f0ef853e,
        64'h45912000_061343dc,
        64'hfd843783_c2e19423,
        64'h474dbf9f_f0ef853e,
        64'h03a00593_460143dc,
        64'hfd843783_c0bff0ef,
        64'h853e0380_05934601,
        64'h43dcfd84_3783c1df,
        64'hf0ef853a_03600593,
        64'h3ff78613_67bd43d8,
        64'hfd843783_c33ff0ef,
        64'h853a0340_0593eff7,
        64'h861367c1_43d8fd84,
        64'h3783cc9f_f0ef853e,
        64'h02800593_464143dc,
        64'hfd843783_cdbff0ef,
        64'h853a0290_0593863e,
        64'h0ff7f793_0017e793,
        64'hfeb44783_43d8fd84,
        64'h3783fe04_05a3a019,
        64'hfef405a3_47a9c789,
        64'h27818ff9_040007b7,
        64'h873e579c_fd843783,
        64'ha005fef4_05a347b1,
        64'hc7892781_8ff90200,
        64'h07b7873e_579cfd84,
        64'h3783a82d_fef405a3,
        64'h47b9c789_27818ff9,
        64'h010007b7_873e579c,
        64'hfd843783_a8c5fef4,
        64'h26234785_c7892781,
        64'hfec42783_fef42623,
        64'h87aa0c00_30effd84,
        64'h3503a807_85930006,
        64'h27b7b19f_f0ef0c80,
        64'h051300f7_16634000,
        64'h07b7873e_27818ff9,
        64'hc00007b7_873e579c,
        64'hfd843783_02f71363,
        64'h4789873e_0367c783,
        64'hfd843783_da3ff0ef,
        64'h853e0290_0593463d,
        64'h43dcfd84_3783a811,
        64'hdb7ff0ef_853e0290,
        64'h0593463d_43dcfd84,
        64'h378300f7_1c634789,
        64'h873e0367_c783fd84,
        64'h3783d798_fd843783,
        64'h0007871b_87aac8ff,
        64'hf0ef853e_93811782,
        64'h27810407_879b43dc,
        64'hfd843783_02e78b23,
        64'hfd843783_0ff7f713,
        64'h87aad4ff_f0ef853e,
        64'h0fe00593_43dcfd84,
        64'h3783f3e5_27818b85,
        64'h2781fea4_4783fef4,
        64'h052387aa_df1ff0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_a821fef4,
        64'h052387aa_e09ff0ef,
        64'h853e02f0_059343dc,
        64'hfd843783_e53ff0ef,
        64'h853e02f0_05934605,
        64'h43dcfd84_3783c0df,
        64'hf0ef3e80_0513e6df,
        64'hf0ef853e_02900593,
        64'h460143dc_fd843783,
        64'ha811e81f_f0ef853e,
        64'h02900593_464143dc,
        64'hfd843783_ac354785,
        64'hc2e1a223_4705a33f,
        64'hf0ef0625_05130000,
        64'h45170625_85930000,
        64'h45970b50_0613a015,
        64'h02f71e63_4789873e,
        64'h27810ff7_f7932781,
        64'h87aae0ff_f0ef853e,
        64'h0fe00593_43dcfd84,
        64'h37830607_b823fd84,
        64'h3783d7f8_4719fd84,
        64'h37830607_a223fd84,
        64'h378302e7_8023fd84,
        64'h37830207_c703fd04,
        64'h3783cfd8_fd843783,
        64'h4fd8fd04_3783cf98,
        64'hfd843783_4f98fd04,
        64'h3783cbd8_fd843783,
        64'h4bd8fd04_3783cb98,
        64'hfd843783_4b98fd04,
        64'h3783c7d8_fd843783,
        64'h47d8fd04_3783d3d8,
        64'h1117071b_11111737,
        64'hfd843783_c798fd84,
        64'h37834798_fd043783,
        64'hc3d8fcc4_2703fd84,
        64'h378300e7_9023fd84,
        64'h37830007_d703fd04,
        64'h3783c201_a223ae39,
        64'h4785c2e1_a2234705,
        64'hb15ff0ef_14450513,
        64'h00004517_14458593,
        64'h00004597_0b400613,
        64'ha015c3fd_fd043783,
        64'hc201a223_c799fd84,
        64'h3783fcf4_262387b2,
        64'hfcb43823_fca43c23,
        64'h0080f822_fc067139,
        64'h80826105_644260e2,
        64'h0001e8df_f0ef853e,
        64'h85bafea4_47039381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef40523_87bafef4,
        64'h05a387b6_fef42623,
        64'h873286ae_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e2853e,
        64'h87aae7ff_f0ef853e,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_05a387ba,
        64'hfef42623_872e87aa,
        64'h1000e822_ec061101,
        64'h80826105_644260e2,
        64'h0001f39f_f0ef853e,
        64'h85bafe84_57039381,
        64'h17822781_9fb9fec4,
        64'h27032781_feb44783,
        64'hfef41423_87bafef4,
        64'h05a387b6_fef42623,
        64'h873286ae_87aa1000,
        64'he822ec06_11018082,
        64'h61056442_60e2853e,
        64'h87aaf1df_f0ef853e,
        64'h93811782_27819fb9,
        64'hfec42703_2781feb4,
        64'h4783fef4_05a387ba,
        64'hfef42623_872e87aa,
        64'h1000e822_ec061101,
        64'h80826145_74220001,
        64'hc398fd44_2703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_2a2387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61457422,
        64'h000100e7_9023fd64,
        64'h5703fe84_3783fef4,
        64'h3423fd84_3783fcf4,
        64'h1b2387ae_fca43c23,
        64'h1800f422_71798082,
        64'h61457422_000100e7,
        64'h8023fd74_4703fe84,
        64'h3783fef4_3423fd84,
        64'h3783fcf4_0ba387ae,
        64'hfca43c23_1800f422,
        64'h71798082_61056462,
        64'h853e2781_439cfe84,
        64'h3783fea4_34231000,
        64'hec221101_80826105,
        64'h6462853e_93c117c2,
        64'h0007d783_fe843783,
        64'hfea43423_1000ec22,
        64'h11018082_61056462,
        64'h853e0ff7_f7930007,
        64'hc783fe84_3783fea4,
        64'h34231000_ec221101,
        64'h80826145_7422853e,
        64'hfe843783_fae7f5e3,
        64'h47850007_871bfe44,
        64'h2783fef4_22232785,
        64'hfe442783_a829fef4,
        64'h342397ba_1ac70713,
        64'h1ffee717_078a97ba,
        64'h078e87ba_fe446703,
        64'h02f71063_27812701,
        64'hfde45703_0007d783,
        64'h97ba1de6_8713078a,
        64'h97ba078e_87bafe44,
        64'h67031ffe_e697a0b9,
        64'hfe042223_fe043423,
        64'hfcf41f23_87aa1800,
        64'hf4227179_80826145,
        64'h740270a2_0001fef7,
        64'h68e3fe04_3783fe84,
        64'h3703fea4_3423fbff,
        64'hf0effef4_302397ba,
        64'hfe843783_873e078a,
        64'h97ba078a_87bafd84,
        64'h3703fea4_3423fdff,
        64'hf0effca4_3c231800,
        64'hf022f406_71798082,
        64'h01416422_853e639c,
        64'h17e10200_c7b70800,
        64'he4221141_80826109,
        64'h640660a6_853efec4,
        64'h2783fef4_262387aa,
        64'hb38ff0ef_c2650513,
        64'hfffff517_85be567d,
        64'hfb843683_fd040793,
        64'hfe043703_fcf43c23,
        64'hfc043783_fcf43823,
        64'hfc843783_fef43023,
        64'hfd878793_03040793,
        64'h03143423_03043023,
        64'hec1ce818_e414fac4,
        64'h3c23fcb4_3023fca4,
        64'h34230880_e0a2e486,
        64'h71198082_61457402,
        64'h70a2853e_87aab9ef,
        64'hf0efbf65_0513ffff,
        64'hf517fe84_3583fe04,
        64'h3603fd84_3683fd04,
        64'h3703fcd4_3823fcc4,
        64'h3c23feb4_3023fea4,
        64'h34231800_f022f406,
        64'h71798082_61457402,
        64'h70a2853e_87aabdef,
        64'hf0efc945_0513ffff,
        64'hf51785be_567dfd84,
        64'h3683fd04_3703fe84,
        64'h0793fcb4_3823fca4,
        64'h3c231800_f022f406,
        64'h71798082_61657442,
        64'h70e2853e_fec42783,
        64'hfef42623_87aac1ef,
        64'hf0efc765_0513ffff,
        64'hf517fd84_3583fd04,
        64'h3603fc84_3683873e,
        64'hfe043783_fef43023,
        64'hfd878793_03040793,
        64'h03143423_03043023,
        64'hec1ce818_e414fcc4,
        64'h3423fcb4_3823fca4,
        64'h3c230080_f822fc06,
        64'h71598082_61257402,
        64'h70a2853e_fec42783,
        64'hfef42623_87aac7ef,
        64'hf0efcd65_0513ffff,
        64'hf517fd84_3583567d,
        64'hfd043683_873efe04,
        64'h3783fef4_3023fd07,
        64'h87930304_07930314,
        64'h34230304_3023ec1c,
        64'he818e414_e010fcb4,
        64'h3823fca4_3c231800,
        64'hf022f406_711d8082,
        64'h61097442_70e2853e,
        64'hfec42783_fef42623,
        64'h87aacdaf_f0efd905,
        64'h0513ffff_f51785be,
        64'h567dfc84_3683fd84,
        64'h0793fe04_3703fef4,
        64'h3023fc87_87930404,
        64'h07930314_3c230304,
        64'h3823f41c_f018ec14,
        64'he810e40c_fca43423,
        64'h0080f822_fc067119,
        64'h8082610d_644a60ea,
        64'h853e2781_fd843783,
        64'h97024501_f9043583,
        64'h863ef884_3683f984,
        64'h3703fd84_3783a019,
        64'h17fdf884_378300f7,
        64'h6663f884_3783fd84,
        64'h3703d807_99630007,
        64'hc783f804_37830001,
        64'hf8f43023_0785f804,
        64'h37839702_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_37830007,
        64'hc503f804_3783a80d,
        64'hf8f43023_0785f804,
        64'h37839702_02500513,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h3783a8b9_f8f43023,
        64'h0785f804_3783fca4,
        64'h3c23ba2f_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_36838736,
        64'h47814841_88bae03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_270386be,
        64'h639cf6e4_3c230087,
        64'h8713f784_3783a089,
        64'hfca43c23_cfcff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h87364781_484188ba,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442703,
        64'h86be639c_f6e43c23,
        64'h00878713_f7843783,
        64'hc3b10ff7_f793fbb4,
        64'h4783faf4_0da34785,
        64'hfef42623_0217e793,
        64'hfec42783_fef42423,
        64'h47c1a239_f8f43023,
        64'h0785f804_3783fce7,
        64'he7e32701_fe842703,
        64'hfce42223_0017871b,
        64'hfc442783_97020200,
        64'h0513f904_3583863e,
        64'hf8843683_f9843703,
        64'hfce43c23_00178713,
        64'hfd843783_a00dcf8d,
        64'h27818b89_fec42783,
        64'hfbcdfee4_2223fff7,
        64'h871bfe44_2783d3e1,
        64'h27814007_f793fec4,
        64'h2783cf91_0007c783,
        64'hfc843783_9702f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'h0007c503_fce43423,
        64'h00178713_fc843783,
        64'ha03dfce7_e7e32701,
        64'hfe842703_fce42223,
        64'h0017871b_fc442783,
        64'h97020200_0513f904,
        64'h3583863e_f8843683,
        64'hf9843703_fce43c23,
        64'h00178713_fd843783,
        64'ha00de7a5_27818b89,
        64'hfec42783_fcf42223,
        64'h87b200d7_73630006,
        64'h071b0007_869bfe44,
        64'h2783fc44_2603cf91,
        64'h27814007_f793fec4,
        64'h2783fcf4_222387aa,
        64'h8aaff0ef_fc843503,
        64'h85be57fd_a011fe44,
        64'h6783c781_2781fe44,
        64'h2783fcf4_3423639c,
        64'hf6e43c23_00878713,
        64'hf7843783_a4a1f8f4,
        64'h30230785_f8043783,
        64'hfce7e7e3_2701fe84,
        64'h2703fce4_28230017,
        64'h871bfd04_27839702,
        64'h02000513_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_3783a00d,
        64'hcf8d2781_8b89fec4,
        64'h27839702_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_37830ff7,
        64'hf513439c_f6e43c23,
        64'h00878713_f7843783,
        64'hfce7e7e3_2701fe84,
        64'h2703fce4_28230017,
        64'h871bfd04_27839702,
        64'h02000513_f9043583,
        64'h863ef884_3683f984,
        64'h3703fce4_3c230017,
        64'h8713fd84_3783a00d,
        64'hef8d2781_8b89fec4,
        64'h2783fcf4_28234785,
        64'ha631f8f4_30230785,
        64'hf8043783_fca43c23,
        64'he50ff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_47818836,
        64'h88b2e03e_fe842783,
        64'he43efec4_2783fe44,
        64'h2603fd44_6683fb44,
        64'h6703faf4_2a232781,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783a801,
        64'h278193c1_17c2439c,
        64'hf6e43c23_00878713,
        64'hf7843783_cf812781,
        64'h0807f793_fec42783,
        64'ha8152781_0ff7f793,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783cf81,
        64'h27810407_f793fec4,
        64'h2783a841_fca43c23,
        64'hee0ff0ef_f9843503,
        64'hf9043583_fd843603,
        64'hf8843683_47818836,
        64'h88b2e03e_fe842783,
        64'he43efec4_2783fe44,
        64'h2603fd44_66836398,
        64'hf6e43c23_00878713,
        64'hf7843783_c3b12781,
        64'h1007f793_fec42783,
        64'ha8f9fca4_3c23847f,
        64'hf0eff984_3503f904,
        64'h3583fd84_3603f884,
        64'h36834781_883688b2,
        64'he03efe84_2783e43e,
        64'hfec42783_fe442603,
        64'hfd446683_6398f6e4,
        64'h3c230087_8713f784,
        64'h3783c3b1_27812007,
        64'hf793fec4_2783a235,
        64'hfca43c23_f7cff0ef,
        64'hf9843503_f9043583,
        64'hfd843603_f8843683,
        64'h87b68832_88aee03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_2583fd44,
        64'h66030ff7_f69301f7,
        64'hd79bfb04_27839301,
        64'h02079713_27812781,
        64'h40f707bb_8f3dfb04,
        64'h270341f7_d79bfb04,
        64'h2783faf4_2823439c,
        64'hf6e43c23_00878713,
        64'hf7843783_a8012781,
        64'h4107d79b_0107979b,
        64'h439cf6e4_3c230087,
        64'h8713f784_3783cf91,
        64'h27810807_f793fec4,
        64'h2783a81d_27810ff7,
        64'hf793439c_f6e43c23,
        64'h00878713_f7843783,
        64'hcf812781_0407f793,
        64'hfec42783_a2cdfca4,
        64'h3c23833f_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_3683872e,
        64'h87ba8836_88b2e03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_2603fd44,
        64'h66830ff7_f71393fd,
        64'hfa843783_85be8f99,
        64'h8fb9fa84_378343f7,
        64'hd713fa84_3783faf4,
        64'h3423639c_f6e43c23,
        64'h00878713_f7843783,
        64'hc3bd2781_1007f793,
        64'hfec42783_ac89fca4,
        64'h3c239bbf_f0eff984,
        64'h3503f904_3583fd84,
        64'h3603f884_3683872e,
        64'h87ba8836_88b2e03e,
        64'hfe842783_e43efec4,
        64'h2783fe44_2603fd44,
        64'h66830ff7_f71393fd,
        64'hfa043783_85be8f99,
        64'h8fb9fa04_378343f7,
        64'hd713fa04_3783faf4,
        64'h3023639c_f6e43c23,
        64'h00878713_f7843783,
        64'hc3bd2781_2007f793,
        64'hfec42783_18f71d63,
        64'h06400793_873e0007,
        64'hc783f804_378300f7,
        64'h0b630690_0793873e,
        64'h0007c783_f8043783,
        64'hfef42623_9bf9fec4,
        64'h2783c791_27814007,
        64'hf793fec4_2783fef4,
        64'h26239bcd_fec42783,
        64'h00f70763_06400793,
        64'h873e0007_c783f804,
        64'h378302f7_00630690,
        64'h0793873e_0007c783,
        64'hf8043783_fef42623,
        64'h0207e793_fec42783,
        64'h00f71863_05800793,
        64'h873e0007_c783f804,
        64'h3783fef4_26239bbd,
        64'hfec42783_fcf42a23,
        64'h47a9a809_fcf42a23,
        64'h478900f7_16630620,
        64'h0793873e_0007c783,
        64'hf8043783_a035fcf4,
        64'h2a2347a1_00f71663,
        64'h06f00793_873e0007,
        64'hc783f804_3783a099,
        64'hfcf42a23_47c100f7,
        64'h16630580_0793873e,
        64'h0007c783_f8043783,
        64'h00f70b63_07800793,
        64'h873e0007_c783f804,
        64'h37838782_97babee7,
        64'h87930000_57970007,
        64'h871b439c_97babfe7,
        64'h87930000_57970027,
        64'h97139381_02069793,
        64'h6ce7e363_05300793,
        64'h0006871b_fdb7869b,
        64'h27810007_c783f804,
        64'h37830001_a0110001,
        64'ha0210001_a031f8f4,
        64'h30230785_f8043783,
        64'hfef42623_1007e793,
        64'hfec42783_a015f8f4,
        64'h30230785_f8043783,
        64'hfef42623_1007e793,
        64'hfec42783_a835f8f4,
        64'h30230785_f8043783,
        64'hfef42623_1007e793,
        64'hfec42783_a889f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0407e793,
        64'hfec42783_06f71663,
        64'h06800793_873e0007,
        64'hc783f804_3783f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0807e793,
        64'hfec42783_a079f8f4,
        64'h30230785_f8043783,
        64'hfef42623_2007e793,
        64'hfec42783_0af71463,
        64'h06c00793_873e0007,
        64'hc783f804_3783f8f4,
        64'h30230785_f8043783,
        64'hfef42623_1007e793,
        64'hfec42783_878297ba,
        64'hcb478793_00005797,
        64'h0007871b_439c97ba,
        64'hcc478793_00005797,
        64'h00279713_93810206,
        64'h97930ee7_e96347c9,
        64'h0006871b_f987869b,
        64'h27810007_c783f804,
        64'h3783f8f4_30230785,
        64'hf8043783_fef42223,
        64'h27814781_00075363,
        64'h0007871b_fbc42783,
        64'hfaf42e23_439cf6e4,
        64'h3c230087_8713f784,
        64'h378302f7_1a6302a0,
        64'h0793873e_0007c783,
        64'hf8043783_a091fef4,
        64'h222387aa_f86ff0ef,
        64'h853ef804_0793cb91,
        64'h87aaf54f_f0ef853e,
        64'h0007c783_f8043783,
        64'hf8f43023_0785f804,
        64'h3783fef4_26234007,
        64'he793fec4_278308f7,
        64'h106302e0_0793873e,
        64'h0007c783_f8043783,
        64'hfe042223_f8f43023,
        64'h0785f804_3783fef4,
        64'h2423fc04_2783a029,
        64'hfef42423_278140f0,
        64'h07bbfc04_2783fef4,
        64'h26230027_e793fec4,
        64'h27830207_d0632781,
        64'hfc042783_fcf42023,
        64'h439cf6e4_3c230087,
        64'h8713f784_378304f7,
        64'h176302a0_0793873e,
        64'h0007c783_f8043783,
        64'ha8b9fef4_242387aa,
        64'h833ff0ef_853ef804,
        64'h0793cb91_87aa801f,
        64'hf0ef853e_0007c783,
        64'hf8043783_fe042423,
        64'hf3852781_fe042783,
        64'h0001fe04_2023a021,
        64'hfef42023_4785f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0107e793,
        64'hfec42783_a01dfef4,
        64'h20234785_f8f43023,
        64'h0785f804_3783fef4,
        64'h26230087_e793fec4,
        64'h2783a091_fef42023,
        64'h4785f8f4_30230785,
        64'hf8043783_fef42623,
        64'h0047e793_fec42783,
        64'ha08dfef4_20234785,
        64'hf8f43023_0785f804,
        64'h3783fef4_26230027,
        64'he793fec4_2783a041,
        64'hfef42023_4785f8f4,
        64'h30230785_f8043783,
        64'hfef42623_0017e793,
        64'hfec42783_878297ba,
        64'he6878793_00005797,
        64'h0007871b_439c97ba,
        64'he7878793_00005797,
        64'h00279713_93810206,
        64'h97930ce7_e06347c1,
        64'h0006871b_fe07869b,
        64'h27810007_c783f804,
        64'h3783fe04_2623f8f4,
        64'h30230785_f8043783,
        64'h2270006f_f8f43023,
        64'h0785f804_37839702,
        64'hf9043583_863ef884,
        64'h3683f984_3703fce4,
        64'h3c230017_8713fd84,
        64'h37830007_c503f804,
        64'h378302f7_0b630250,
        64'h0793873e_0007c783,
        64'hf8043783_26b0006f,
        64'hf8f43c23_86678793,
        64'h00000797_26079de3,
        64'hf9043783_fc043c23,
        64'hf6e43c23_f8d43023,
        64'hf8c43423_f8b43823,
        64'hf8a43c23_1100e922,
        64'hed067135_8082610d,
        64'h644a60ea_853e87aa,
        64'hb47ff0ef_fb843503,
        64'hfb043583_fa843603,
        64'hfa043683_fe843783,
        64'h883688b2_e03ef904,
        64'h2783e43e_401ce83e,
        64'h441cfc04_0713f974,
        64'h46830007_861bf884,
        64'h3783f6e7_ffe347fd,
        64'hfe843703_c791f984,
        64'h3783f8f4_3c2302f7,
        64'h57b3f884_3783f984,
        64'h3703fcf7_08239736,
        64'hff040693_fed43423,
        64'h00170693_fe843703,
        64'h0ff7f793_37d90ff7,
        64'hf7939fb9_fe744703,
        64'h06100793_a0190410,
        64'h0793c781_27810207,
        64'hf793441c_a01d0ff7,
        64'hf7930307_879bfe74,
        64'h478300e7_e96347a5,
        64'h0ff7f713_fe744783,
        64'hfef403a3_02f777b3,
        64'hf8843783_f9843703,
        64'hc7c1f984_3783c781,
        64'h27814007_f793441c,
        64'hc41c9bbd_441ce781,
        64'hf9843783_fe043423,
        64'hf8f42823_87baf8f4,
        64'h0ba38746_f9043423,
        64'hf8e43c23_fad43023,
        64'hfac43423_fab43823,
        64'hfaa43c23_1100e922,
        64'hed067135_8082610d,
        64'h644a60ea_853e87aa,
        64'hc5fff0ef_fb843503,
        64'hfb043583_fa843603,
        64'hfa043683_fe843783,
        64'h883688b2_e03ef904,
        64'h2783e43e_401ce83e,
        64'h441cfc04_0713f974,
        64'h46830007_861bf884,
        64'h3783f6e7_ffe347fd,
        64'hfe843703_c791f984,
        64'h3783f8f4_3c2302f7,
        64'h57b3f884_3783f984,
        64'h3703fcf7_08239736,
        64'hff040693_fed43423,
        64'h00170693_fe843703,
        64'h0ff7f793_37d90ff7,
        64'hf7939fb9_fe744703,
        64'h06100793_a0190410,
        64'h0793c781_27810207,
        64'hf793441c_a01d0ff7,
        64'hf7930307_879bfe74,
        64'h478300e7_e96347a5,
        64'h0ff7f713_fe744783,
        64'hfef403a3_02f777b3,
        64'hf8843783_f9843703,
        64'hc7c1f984_3783c781,
        64'h27814007_f793441c,
        64'hc41c9bbd_441ce781,
        64'hf9843783_fe043423,
        64'hf8f42823_87baf8f4,
        64'h0ba38746_f9043423,
        64'hf8e43c23_fad43023,
        64'hfac43423_fab43823,
        64'hfaa43c23_1100e922,
        64'hed067135_80826161,
        64'h640660a6_853e87aa,
        64'hc65ff0ef_fe843503,
        64'hfe043583_fd843603,
        64'hfd043683_fc843703,
        64'hfc043783_883e88ba,
        64'h441c4818_00e78023,
        64'h02000713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_3783cf91,
        64'h27818ba1_481ca015,
        64'h00e78023_02b00713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h3783cf99_27818b91,
        64'h481ca0a1_00e78023,
        64'h02d00713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_3783cf99,
        64'h0ff7f793_fbf44783,
        64'h06e7e863_47fdfc04,
        64'h370300e7_80230300,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_00e7ef63,
        64'h47fdfc04_370300e7,
        64'h80230620_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'h00e7ef63_47fdfc04,
        64'h370302f7_14634789,
        64'h0007871b_fb842783,
        64'ha81500e7_80230580,
        64'h071397ba_fc843703,
        64'hfce43023_00178713,
        64'hfc043783_02e7e063,
        64'h47fdfc04_3703c785,
        64'h27810207_f793481c,
        64'h02f71a63_47c10007,
        64'h871bfb84_2783a88d,
        64'h00e78023_07800713,
        64'h97bafc84_3703fce4,
        64'h30230017_8713fc04,
        64'h378302e7_e06347fd,
        64'hfc043703_e7852781,
        64'h0207f793_481c02f7,
        64'h1a6347c1_0007871b,
        64'hfb842783_fcf43023,
        64'h17fdfc04_378300f7,
        64'h176347c1_0007871b,
        64'hfb842783_cf89fc04,
        64'h3783fcf4_302317fd,
        64'hfc043783_02f71663,
        64'hfc043703_00846783,
        64'h00f70863_fc043703,
        64'h00046783_c3a9fc04,
        64'h3783e7a1_27814007,
        64'hf793481c_12078363,
        64'h27818bc1_481cfce7,
        64'hf6e347fd_fc043703,
        64'h00f77763_fc043703,
        64'h00846783_cf812781,
        64'h8b85481c_00e78023,
        64'h03000713_97bafc84,
        64'h3703fce4_30230017,
        64'h8713fc04_3783a831,
        64'hfce7fae3_47fdfc04,
        64'h370302f7_7563fc04,
        64'h37030004_678300e7,
        64'h80230300_071397ba,
        64'hfc843703_fce43023,
        64'h00178713_fc043783,
        64'ha831c41c_37fd441c,
        64'hc3952781_8bb1481c,
        64'he7890ff7_f793fbf4,
        64'h4783cb9d_27818b85,
        64'h481ccf9d_2781441c,
        64'hebd12781_8b89481c,
        64'hfaf42c23_87bafaf4,
        64'h0fa38746_87c2fcf4,
        64'h3023fce4_3423fcd4,
        64'h3823fcc4_3c23feb4,
        64'h3023fea4_34230880,
        64'he0a2e486_715d8082,
        64'h61256446_60e6853e,
        64'hfc843783_fcf769e3,
        64'hfac46783_8f1dfe04,
        64'h3783fc84_37039702,
        64'h02000513_fd043583,
        64'h863efc04_3683fd84,
        64'h3703fce4_34230017,
        64'h8713fc84_3783a00d,
        64'hcb9d2781_8b89fa84,
        64'h2783f7e1_fb043783,
        64'h9702fd04_3583863e,
        64'hfc043683_fd843703,
        64'hfce43423_00178713,
        64'hfc843783_0007c503,
        64'h97bafb04_3783fb84,
        64'h3703faf4_382317fd,
        64'hfb043783_a81dfcf7,
        64'h67e3fe84_3703fac4,
        64'h6783fef4_34230785,
        64'hfe843783_97020200,
        64'h0513fd04_3583863e,
        64'hfc043683_fd843703,
        64'hfce43423_00178713,
        64'hfc843783_a035fef4,
        64'h3423fb04_3783efa5,
        64'h27818b85_fa842783,
        64'he3c92781_8b89fa84,
        64'h2783fef4_3023fc84,
        64'h3783faf4_242387ba,
        64'hfaf42623_874687c2,
        64'hfaf43823_fae43c23,
        64'hfcd43023_fcc43423,
        64'hfcb43823_fca43c23,
        64'h1080e8a2_ec86711d,
        64'h80826145_740270a2,
        64'h853efec4_2783ffc5,
        64'h87aaf6df_f0ef853e,
        64'h0007c783_639cfd84,
        64'h3783fef4_2623fd07,
        64'h879b2781_9fb92781,
        64'h0007c783_e290fd84,
        64'h36830017_8613639c,
        64'hfd843783_0007871b,
        64'h0017979b_9fb90027,
        64'h979b87ba_fec42703,
        64'ha825fe04_2623fca4,
        64'h3c231800_f022f406,
        64'h71798082_61056462,
        64'h853e0ff7_f7938b85,
        64'h4781a011_478500e7,
        64'he4630390_07930ff7,
        64'hf713fef4_478300e7,
        64'hfc6302f0_07930ff7,
        64'hf713fef4_4783fef4,
        64'h07a387aa_1000ec22,
        64'h11018082_61457422,
        64'h853e2781_40f707b3,
        64'hfd843783_fe843703,
        64'hf3e5fce4_3823fff7,
        64'h8713fd04_3783cb81,
        64'h0007c783_fe843783,
        64'hfef43423_0785fe84,
        64'h3783a031_fef43423,
        64'hfd843783_fcb43823,
        64'hfca43c23_1800f422,
        64'h71798082_61457402,
        64'h70a20001_9682853e,
        64'h85bafef4_47836798,
        64'hfe043783_6394fe04,
        64'h3783cf81_0ff7f793,
        64'hfef44783_fef407a3,
        64'hfcd43823_fcc43c23,
        64'hfeb43023_87aa1800,
        64'hf022f406_71798082,
        64'h61457402_70a20001,
        64'h8e7ff0ef_853efef4,
        64'h4783c791_0ff7f793,
        64'hfef44783_fef407a3,
        64'hfcd43823_fcc43c23,
        64'hfeb43023_87aa1800,
        64'hf022f406_71798082,
        64'h61457422_0001fef4,
        64'h07a3fcd4_3823fcc4,
        64'h3c23feb4_302387aa,
        64'h1800f422_71798082,
        64'h61457422_000100e7,
        64'h8023fef4_470397ba,
        64'hfd843783_fe043703,
        64'h00f77b63_fd043783,
        64'hfd843703_fef407a3,
        64'hfcd43823_fcc43c23,
        64'hfeb43023_87aa1800,
        64'hf4227179_8082610d,
        64'h690a64aa_644a60ea,
        64'hf6040113_853e8126,
        64'h814a4781_2b0010ef,
        64'h6f050513_00005517,
        64'ha80157f9_2c0010ef,
        64'h4b050513_00005517,
        64'h85befac4_27832d20,
        64'h10ef4aa5_05130000,
        64'h5517c395_2781fac4,
        64'h2783faf4_262387aa,
        64'hb63ff0ef_f6843503,
        64'h85be863a_f6442703,
        64'h2781739c_f8043783,
        64'h304010ef_72c50513,
        64'h00005517_f8f43023,
        64'hf8843783_eae7d2e3,
        64'h478d0007_871bfd04,
        64'h2783fcf4_28232785,
        64'hfd042783_330010ef,
        64'h57850513_00005517,
        64'hfce7d6e3_04700793,
        64'h0007871b_fdc42783,
        64'hfcf42e23_2785fdc4,
        64'h27833560_10ef6f65,
        64'h05130000_551785be,
        64'h27810387_c78397ba,
        64'hfdc42783_f7843703,
        64'ha02dfc04_2e2337a0,
        64'h10ef78a5_05130000,
        64'h55173860_10ef77e5,
        64'h05130000_551785be,
        64'h7b9cf784_378339a0,
        64'h10ef77a5_05130000,
        64'h551785be_779cf784,
        64'h37833ae0_10ef7765,
        64'h05130000_551785be,
        64'h739cf784_3783fce7,
        64'hd7e347bd_0007871b,
        64'hfd842783_fcf42c23,
        64'h2785fd84_27833da0,
        64'h10ef77a5_05130000,
        64'h551785be_27810107,
        64'hc78397ba_fd842783,
        64'hf7843703_a02dfc04,
        64'h2c233fe0_10ef7a65,
        64'h05130000_5517fce7,
        64'hd7e347bd_0007871b,
        64'hfd442783_fcf42a23,
        64'h2785fd44_27834220,
        64'h10ef7c25_05130000,
        64'h551785be_27810007,
        64'hc78397ba_fd442783,
        64'hf7843703_a02dfc04,
        64'h2a234460_10ef7c65,
        64'h05130000_55174520,
        64'h10ef7ba5_05130000,
        64'h551785be_fd042783,
        64'hf6f43c23_97ba2701,
        64'h0077171b_fd042703,
        64'hf8843783_aa91fc04,
        64'h2823aac9_57f94820,
        64'h10ef7ca5_05130000,
        64'h551785be_fac42783,
        64'h494010ef_66c50513,
        64'h00005517_c3952781,
        64'hfac42783_faf42623,
        64'h87aad25f_f0ef853a,
        64'h85be4605_278167bc,
        64'hfa043783_f8843703,
        64'hf8f43423_00078793,
        64'h878a40f1_01330792,
        64'h839107bd_f8e43823,
        64'h177d873e_893a870a,
        64'hfc043783_4e8010ef,
        64'h81050513_00006517,
        64'h85be4bfc_fa043783,
        64'h4fc010ef_80450513,
        64'h00006517_85be4bbc,
        64'hfa043783_510010ef,
        64'h7f050513_00005517,
        64'h85be67bc_fa043783,
        64'h524010ef_7ec50513,
        64'h00005517_85be739c,
        64'hfa043783_538010ef,
        64'h7e850513_00005517,
        64'h85be6f9c_fa043783,
        64'h54c010ef_7e450513,
        64'h00005517_85be4bdc,
        64'hfa043783_560010ef,
        64'h7e050513_00005517,
        64'h85be4b9c_fa043783,
        64'h574010ef_7dc50513,
        64'h00005517_85be47dc,
        64'hfa043783_588010ef,
        64'h7d850513_00005517,
        64'h85be479c_fa043783,
        64'h59c010ef_7e450513,
        64'h00005517_fce7d7e3,
        64'h479d0007_871bfcc4,
        64'h2783fcf4_26232785,
        64'hfcc42783_5c0010ef,
        64'h80050513_00006517,
        64'h85be2781_0007c783,
        64'h97baf984_3703fcc4,
        64'h2783a02d_fc042623,
        64'hf8f43c23_fa043783,
        64'h5ec010ef_81c50513,
        64'h00006517_5f8010ef,
        64'h80850513_00006517,
        64'hfaf43023_fb043783,
        64'ha68d57f9_610010ef,
        64'h80050513_00006517,
        64'h85befac4_27836220,
        64'h10ef7fa5_05130000,
        64'h5517c395_2781fac4,
        64'h2783faf4_262387aa,
        64'heb3ff0ef_853e4585,
        64'h4605fb04_3783faf4,
        64'h38230007_8793878a,
        64'h40f10133_07928391,
        64'h07bdfae4_3c23177d,
        64'h873efc04_3783fcf4,
        64'h30232000_07936720,
        64'h10ef8325_05130000,
        64'h6517aed1_57fd6820,
        64'h10ef81a5_05130000,
        64'h6517cb89_2781fc84,
        64'h2783fcf4_242387aa,
        64'he5bff0ef_84be878a,
        64'hf6f42223_87aef6a4,
        64'h34231100_e14ae526,
        64'he922ed06_71358082,
        64'h61457402_70a2853e,
        64'h4781a011_57fd6ca0,
        64'h10ef8425_05130000,
        64'h651785be_fe442783,
        64'hcf812781_fe442783,
        64'hfef42223_87aa7600,
        64'h30efc2a5_05131fff,
        64'h051785be_863afe84,
        64'h3683fd44_2783fd04,
        64'h2703fae7_e0e3678d,
        64'h0007871b_fd042783,
        64'hfef43423_97ba0060,
        64'h07b7fe84_3703fcf4,
        64'h28239fb9_77f5fd04,
        64'h2703a0b5_57fd7320,
        64'h10ef8aa5_05130000,
        64'h651785be_fe042783,
        64'hcf812781_fe042783,
        64'hfef42023_87aa7c80,
        64'h30efc925_05131fff,
        64'h051785be_660dfe84,
        64'h3683fd44_2783a8a1,
        64'hfef43423_fd843783,
        64'hfcf42823_87bafcf4,
        64'h2a238732_87aefca4,
        64'h3c231800_f022f406,
        64'h71798082_61056442,
        64'h60e2853e_478179a0,
        64'h10ef8f25_05130000,
        64'h6517a801_57f57aa0,
        64'h10ef8d25_05130000,
        64'h651785be_fe442783,
        64'hcf812781_fe442783,
        64'hfef42223_87aa53c0,
        64'h20efd0a5_05131fff,
        64'h0517a081_57f97da0,
        64'h10ef8da5_05130000,
        64'h651785be_fe442783,
        64'hcf812781_fe442783,
        64'hfef42223_87aa4ab0,
        64'h10efd3a5_05131fff,
        64'h0517fe84_3583863e,
        64'h43dcfe84_3783a8b5,
        64'h57fd0170_10ef8f65,
        64'h05130000_6517eb89,
        64'hfe843783_fea43423,
        64'h289010ef_45010330,
        64'h10ef8fa5_05130000,
        64'h65171000_e822ec06,
        64'h11018082_61457402,
        64'h70a20001_eb9ff0ef,
        64'h01078513_07fa478d,
        64'h02000593_ec9ff0ef,
        64'h00878513_07fa478d,
        64'h0c700593_ed9ff0ef,
        64'h00c78513_07fa478d,
        64'h458dee7f_f0ef0047,
        64'h851307fa_478d85be,
        64'h0ff7f793_27810087,
        64'hd79bfec4_2783f03f,
        64'hf0ef01e7_9513478d,
        64'h85be0ff7_f793fec4,
        64'h2783f17f_f0ef00c7,
        64'h851307fa_478d0800,
        64'h0593f27f_f0ef0047,
        64'h851307fa_478d4581,
        64'hfef42623_02f757bb,
        64'hfdc42703_27810047,
        64'h979bfd84_2783fcf4,
        64'h2c2387ba_fcf42e23,
        64'h872e87aa_1800f022,
        64'hf4067179_80826105,
        64'h644260e2_0001f6bf,
        64'hf0ef01e7_9513478d,
        64'h85befef4_4783dfed,
        64'h87aafc9f_f0ef0001,
        64'hfef407a3_87aa1000,
        64'he822ec06_11018082,
        64'h01416402_60a2853e,
        64'h27810207_f7932781,
        64'h87aafd3f_f0ef0147,
        64'h851307fa_478d0800,
        64'he022e406_11418082,
        64'h61056462_853e0ff7,
        64'hf7930007_c783fe84,
        64'h3783fea4_34231000,
        64'hec221101_80826145,
        64'h74220001_00e78023,
        64'hfd744703_fe843783,
        64'hfef43423_fd843783,
        64'hfcf40ba3_87aefca4,
        64'h3c231800_f4227179,
        64'ha00119f0_10efa3e5,
        64'h05130000_65178402,
        64'h00858593_00006597,
        64'h10000437_eb812781,
        64'hfe442783_1c1010ef,
        64'ha3850513_00006517,
        64'hfce7d7e3_47bd0007,
        64'h871bfe84_2783fef4,
        64'h24232785_fe842783,
        64'h1e5010ef_a7c50513,
        64'h00006517_85be2781,
        64'h0007c783_97bafd84,
        64'h3703fe84_2783a02d,
        64'hfe042423_209010ef,
        64'ha8850513_00006517,
        64'h100005b7_fcf43c23,
        64'h100007b7_fef42223,
        64'h87aa3700_00ef1000,
        64'h053765a1_231010ef,
        64'haa850513_00006517,
        64'hfae7d0e3_47890007,
        64'h871bfec4_2783fef4,
        64'h26232785_fec42783,
        64'h255010ef_ac450513,
        64'h00006517_85b6863e,
        64'h43dc97ba_078eeaa7,
        64'h0713fec4_27831fff,
        64'h07174394_97baebc7,
        64'h8793070e_fec42703,
        64'h1fff0797_289010ef,
        64'haf050513_00006517,
        64'h4a7010ef_24078513,
        64'h000f47b7_a8a1fe04,
        64'h26232a70_10efae65,
        64'h05130000_65171be0,
        64'h00efa007_85130262,
        64'h67b72007_859367f1,
        64'h1800f022_f4067179,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_100004b7,
        64'h15058593_00006597,
        64'hf1402573_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_090000ef,
        64'hf9810113_3fff0117,
        64'hfeb56ce3_00450513,
        64'h00052023_00b57863,
        64'hc2a18593_01450513,
        64'h1fff0517_fec5e8e3,
        64'h00458593_00450513,
        64'h0055a023_00052283,
        64'h00c5fc63_03460613,
        64'h1fff0617_fdc58593,
        64'h1fff0597_de450513,
        64'h00007517_84c18193,
        64'h1fff1197_09249063,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
